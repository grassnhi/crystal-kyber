`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/12/2025 01:24:05 PM
// Design Name: 
// Module Name: tb_test_kyber
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module test_kyber_tb;

    // Inputs
    reg clk;
    reg rst;
    reg start;
    reg [1:0] mode;
    reg [255:0] random_coin;
    reg [255:0] m_in;
    reg [6399:0] pk_in;
    reg [6143:0] sk_in;
    reg [6143:0] c_in;

    // Outputs
    wire [255:0] m_out;
    wire [6399:0] pk_out;
    wire [6143:0] sk_out;
    wire [6143:0] c_out;
    wire finish;

    // Instantiate the DUT
    test_kyber uut (
        .clk(clk),
        .rst(rst),
        .start(start),
        .mode(mode),
        .random_coin(random_coin),
        .m_in(m_in),
        .pk_in(pk_in),
        .sk_in(sk_in),
        .c_in(c_in),
        .m_out(m_out),
        .pk_out(pk_out),
        .sk_out(sk_out),
        .c_out(c_out),
        .finish(finish)
    );

    // Clock generation
    initial clk = 0;
    always #5 clk = ~clk; // 100 MHz clock

    initial begin
        // Initialize all inputs
        rst = 1;
        start = 0;
        mode = 0;
        random_coin = 15;
        m_in = 256'hA5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5A5;
        pk_in = 6400'ha4449c1f6511c07619ada306a1498a233a419aa003a305d726a90328209e18da2fc04b4549f6404d535c8b7697c5c7339cdbcb52844cbd338933026f9ecc789c79553141d06d483d579bbc115199b6185f812a08b3a7ae6ef2e26c5763370c5865abfeb6f3b3a9fb18b3736200d22836023b6fd83e74e68302d007c2b125ba3bb814f37f9da65e12f3f60ccb72918b424b66f40768859ca24e060b2e9cb80c43788e5be8307d34bdc375f107b98039fae257e8293a89401ee6d74c91b232a015adf108b8d5537051ef55ab5a5c65a2359a548e77ea6ae7696d91f306dcb69f5b699ce778ae7504c0825f3e791eb4c8c994ea9b027ab79f5caa12117bac01e4598517286616bf572aa284826954f600648c9d15750230a29261d1be519f4daca097fb189a49cd75a71c9a13448b55ab155953a2c68b10a1435cb1a70131f21798b1c2e31772d7fc2ce67ea9f6e16e180812a9d951229367377b7c3bc17ce80f94f7424d839a17f5e57731830a18dc8d022287167f3932f743ca796099c678bae220cb18bbd5027d348506faf19f04c1bfa4ca99f5688b8254484aa46a88b87376dd0d80b097a6b51f446484bcf15c4b8f5cf9e0429978b0c4a877d041549c386d1a2c46c92942c89567a8a3a141248ad0a69aab278d06f95ce4c70cb235cd604798471c2799e47a20438375514bd89c46e0182af6117561dd90113909835656573e58d2a7aae139a2f1b47f4c435457918170c8923575b6599f0eab3e90619b867aee03d0c35e70c778768c08665cbc62ab42d7accdfb303bdc01afc83cb1b64d9383f40952d892db92a15a74744a453885ee2f6176a35c410eaa3acec66a02c07b1624370c1750cd054ac9f72b75306e4bdc63940883bddbce90f3b358fb9995fa77bfe5ce1a2bd6c9e98735733e663594c3cb4d7fc35d61605ebf17293d0ac12780f52d3aec739a8e010598c192d46989aa7320ca0dc15f74858ab8c1530da3d96968308529a50a886174b4397bd92d508c4c1099d9a71a9ebeb5521ff8f7aa30f1295c1989426b28b39f8b4ac442c626160cda08f4026f2b7a49ac130b32fdf598f29e514835c82200bea92b0b72f793c0e5e147b8f2eb9f7a89b0f6945b25;
        sk_in = 6144'hb11bc95746c38e92f249428e35b833ab3031bae51f742958a8513399732c6fb6361e875bcbba030863792f04878f47ebbb97940439241f60414586ba4958b660454013c2a7cf11117e808cb6449e878bf00a26be3c324b7b5a73b96aeabd243a2fe91b652082020a4a04a8dc23281e1016498489323144ef96778680675d4bac0c224467c712a7b3c2ad09d246c309d359dc9cceb42a74a4e88cf19132c63875407f93face116021bf428f5403b24c4ad259c7353629a2083758c977b42140f8b9d19386e347176a0dcfeaa21822a075645ca942fa5a972c598ba075d9da7fa6e04bcc873c86029d55a53d32cc481a4b54ac8350348d83eb6e702910225245859abe6c8672bbcc591f05442e8645a0290eb81b9fc7c80cc121e3787aad9891c8b2e7afbf5afa8414adc827cb196aa8bdb6d37b014fa46562479712860c864bdab8bb81bbcbf42d9a3c32397120a98371b8abca7ba8aa2310d01c9c754b916f6fa6e1952b6e4fe788b7999916dbe64ac12ca3b84578f7af77a2360d520aad27195bb9fd64290bc947a05606858e8ad1a6b52911309e9b68b41844341c065249946e59423b5ff847304a627b018273dbd9327a8f9da0d5667c5716444c1255c893f07a8868487ff78e1c6708c85b9442129eb968f22a5133bca708438291674bb74bbbbd5f902aca85e76a688232d6a61165de699b8a58d0467d78cdab6ad25bf95b3e6a125826ee6572386dd7428e61fa2619b39b6976476ab6cddc79ad8359231a9dc34c20b7a25235fbefa229ce89b65712d9995adca806173a9af8e85e19022dd51b1ffbfb6d92ce6da142bdfcea5408fd75764a74b7de4fa5c13db25a0cfa3a3e41e40d91edc4f8975ef77507d0cc2420798cc97b123aca584c63ba718b3ce3b69e7c5b39d0911ba9a7ac3655c5b7f829fb10071bdd692a59204214ac5b983764fb3b75ab74543cb3c1051b234722b38f3a4ae20af412b960c30c836426808bbfccce9b86d437b6135bd21076aa5089a035b4117c7c03c846282008c4454f6787bbc40a8b06b5698ba0b6dc72301be10de7721df3c759fc261ff3e91177c0;
        c_in = 6144'h2e857cf3867ae53292e5f86f9860041be3dc1db11db66ce377960e79b37f7409a77cb7b58ed3ca7427374f702282d390d1054f58bb8c8402115068bdeaf567b2f4f6dfcac78221c1654b16580ed2f09a0fd601ff826866b155f809ddf0a17bbb04d0bbf0f01efb3379f5471ca19ece5a9844c6086da4d54c5aff31351f06a45346990688c5a775397daad7ad38d3afc961da72cf53559de5476d47a6b2e0e700151bf1340985f2e6f2c60287f8517815b915864998b7227c025d416507d0d430a3d2d57b9b0e064168c52a44e86b84db1a556a9702ddfcdae517f6ef1a9db6c472dd4546cca629e6b3d970f1b5ab468e7240a088c65d8a2cc23f3ef676e7d6f60eb2dd88315fbeacea1cfca380d9ff3d424117842049aa96677467e2092c388ea92e056a37c7eafa10525c6432c957f73ccfafc2c1890268228cfb94c62864329666cf6f713c978b8b92b8867aa6ab5ecaa84526d6bcdba995785a6ebc18c120b2f91faefec247e7a890a8ac8ffd5f2041c09ce73302e239b0e3d50b13fe42cdb70e45fe66d9ad0c508ec72385c284a708446d84af144feb6d4b600bf7ad4921047c8e8dbd6af31756143a5895c2917e3107dcf743294086c3e3da9a3338028047d79d84c6e551670ecf704a4d1977cbd6d1344297f7a5985e8c6203d1e7c0fbf8286fc2a88e84e6baa9556ce7e9be05119a96f34707dd164118c8bd89831e03a142f9f2b441e1675934fbbb2cf8b1608ca010246263eb92b7d3fbff6feb2f350a3462ba02fa56912e768e60a65f399267b8cc2b7a0400f0913da3cffeb4e2699810379b1897e236b606ec668c7b126cbce5f9b3da86d4f8df036f34cf83319cbb486dd6e6329988b50d38db43644d45dee65a13f63745275275f0e8543280d639857c265ec38b06c7578bb493faf01e3b5f49f141c66de49807bbb47d30e7685b9a073673e73f66b69b684f4132c6aa98e5a055754dd6f90423cce4f6a1e075bd4ce9ecb38e0b9299c98a225a0853257f7feebff9af5aa7a9342493b8b115855492371e34757c3c6b49c2e5745df84426151be0c991b0094d93bca8660259ed;

        #100 rst = 0; // Deassert reset

        // --- Mode 0 ---
        #10 mode = 2'd0;
        start = 1;
        #10 start = 0;

        #20 $display("Mode 0:");
        $display("pk_out = %h", pk_out);
        $display("sk_out = %h", sk_out);
        $display("finish = %b", finish);

        // --- Mode 1 ---
        #30 mode = 2'd1;
        start = 1;
        #10 start = 0;

        #20 $display("Mode 1:");
        $display("c_out = %h", c_out);
        $display("finish = %b", finish);

        // --- Mode 2 ---
        #30 mode = 2'd2;
        start = 1;
        #10 start = 0;

        #20 $display("Mode 2:");
        $display("m_out = %h", m_out);
        $display("finish = %b", finish);

        #50;
        $finish;
    end

endmodule

