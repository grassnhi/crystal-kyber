module kcck_round(
    input [1599:0] S_in,        // Input: 5x5 state matrix (1600 bits)
    input wire [4:0] round_index,          // Input: round index (0-23)
    output [1599:0] S_out     // Output: modified 5x5 state matrix
);

    // Intermediate arrays
   wire [63:0] C          [4:0];
   wire [63:0] D          [4:0];
   wire [63:0] A          [4:0][4:0];
   wire [63:0] A_theta    [4:0][4:0];
   wire [63:0] A_rho      [4:0][4:0];
   wire [63:0] A_pi       [4:0][4:0];
   wire [63:0] A_chi      [4:0][4:0];
   reg  [63:0] A_iota     [4:0][4:0];

    // Flatten S_in into 3D array
   assign A[0][0][0]    = S_in[0];
   assign A[1][0][0]    = S_in[64];
   assign A[2][0][0]    = S_in[128];
   assign A[3][0][0]    = S_in[192];
   assign A[4][0][0]    = S_in[256];
   assign A[0][1][0]    = S_in[320];
   assign A[1][1][0]    = S_in[384];
   assign A[2][1][0]    = S_in[448];
   assign A[3][1][0]    = S_in[512];
   assign A[4][1][0]    = S_in[576];
   assign A[0][2][0]    = S_in[640];
   assign A[1][2][0]    = S_in[704];
   assign A[2][2][0]    = S_in[768];
   assign A[3][2][0]    = S_in[832];
   assign A[4][2][0]    = S_in[896];
   assign A[0][3][0]    = S_in[960];
   assign A[1][3][0]    = S_in[1024];
   assign A[2][3][0]    = S_in[1088];
   assign A[3][3][0]    = S_in[1152];
   assign A[4][3][0]    = S_in[1216];
   assign A[0][4][0]    = S_in[1280];
   assign A[1][4][0]    = S_in[1344];
   assign A[2][4][0]    = S_in[1408];
   assign A[3][4][0]    = S_in[1472];
   assign A[4][4][0]    = S_in[1536];
   assign A[0][0][1]    = S_in[1];
   assign A[1][0][1]    = S_in[65];
   assign A[2][0][1]    = S_in[129];
   assign A[3][0][1]    = S_in[193];
   assign A[4][0][1]    = S_in[257];
   assign A[0][1][1]    = S_in[321];
   assign A[1][1][1]    = S_in[385];
   assign A[2][1][1]    = S_in[449];
   assign A[3][1][1]    = S_in[513];
   assign A[4][1][1]    = S_in[577];
   assign A[0][2][1]    = S_in[641];
   assign A[1][2][1]    = S_in[705];
   assign A[2][2][1]    = S_in[769];
   assign A[3][2][1]    = S_in[833];
   assign A[4][2][1]    = S_in[897];
   assign A[0][3][1]    = S_in[961];
   assign A[1][3][1]    = S_in[1025];
   assign A[2][3][1]    = S_in[1089];
   assign A[3][3][1]    = S_in[1153];
   assign A[4][3][1]    = S_in[1217];
   assign A[0][4][1]    = S_in[1281];
   assign A[1][4][1]    = S_in[1345];
   assign A[2][4][1]    = S_in[1409];
   assign A[3][4][1]    = S_in[1473];
   assign A[4][4][1]    = S_in[1537];
   assign A[0][0][2]    = S_in[2];
   assign A[1][0][2]    = S_in[66];
   assign A[2][0][2]    = S_in[130];
   assign A[3][0][2]    = S_in[194];
   assign A[4][0][2]    = S_in[258];
   assign A[0][1][2]    = S_in[322];
   assign A[1][1][2]    = S_in[386];
   assign A[2][1][2]    = S_in[450];
   assign A[3][1][2]    = S_in[514];
   assign A[4][1][2]    = S_in[578];
   assign A[0][2][2]    = S_in[642];
   assign A[1][2][2]    = S_in[706];
   assign A[2][2][2]    = S_in[770];
   assign A[3][2][2]    = S_in[834];
   assign A[4][2][2]    = S_in[898];
   assign A[0][3][2]    = S_in[962];
   assign A[1][3][2]    = S_in[1026];
   assign A[2][3][2]    = S_in[1090];
   assign A[3][3][2]    = S_in[1154];
   assign A[4][3][2]    = S_in[1218];
   assign A[0][4][2]    = S_in[1282];
   assign A[1][4][2]    = S_in[1346];
   assign A[2][4][2]    = S_in[1410];
   assign A[3][4][2]    = S_in[1474];
   assign A[4][4][2]    = S_in[1538];
   assign A[0][0][3]    = S_in[3];
   assign A[1][0][3]    = S_in[67];
   assign A[2][0][3]    = S_in[131];
   assign A[3][0][3]    = S_in[195];
   assign A[4][0][3]    = S_in[259];
   assign A[0][1][3]    = S_in[323];
   assign A[1][1][3]    = S_in[387];
   assign A[2][1][3]    = S_in[451];
   assign A[3][1][3]    = S_in[515];
   assign A[4][1][3]    = S_in[579];
   assign A[0][2][3]    = S_in[643];
   assign A[1][2][3]    = S_in[707];
   assign A[2][2][3]    = S_in[771];
   assign A[3][2][3]    = S_in[835];
   assign A[4][2][3]    = S_in[899];
   assign A[0][3][3]    = S_in[963];
   assign A[1][3][3]    = S_in[1027];
   assign A[2][3][3]    = S_in[1091];
   assign A[3][3][3]    = S_in[1155];
   assign A[4][3][3]    = S_in[1219];
   assign A[0][4][3]    = S_in[1283];
   assign A[1][4][3]    = S_in[1347];
   assign A[2][4][3]    = S_in[1411];
   assign A[3][4][3]    = S_in[1475];
   assign A[4][4][3]    = S_in[1539];
   assign A[0][0][4]    = S_in[4];
   assign A[1][0][4]    = S_in[68];
   assign A[2][0][4]    = S_in[132];
   assign A[3][0][4]    = S_in[196];
   assign A[4][0][4]    = S_in[260];
   assign A[0][1][4]    = S_in[324];
   assign A[1][1][4]    = S_in[388];
   assign A[2][1][4]    = S_in[452];
   assign A[3][1][4]    = S_in[516];
   assign A[4][1][4]    = S_in[580];
   assign A[0][2][4]    = S_in[644];
   assign A[1][2][4]    = S_in[708];
   assign A[2][2][4]    = S_in[772];
   assign A[3][2][4]    = S_in[836];
   assign A[4][2][4]    = S_in[900];
   assign A[0][3][4]    = S_in[964];
   assign A[1][3][4]    = S_in[1028];
   assign A[2][3][4]    = S_in[1092];
   assign A[3][3][4]    = S_in[1156];
   assign A[4][3][4]    = S_in[1220];
   assign A[0][4][4]    = S_in[1284];
   assign A[1][4][4]    = S_in[1348];
   assign A[2][4][4]    = S_in[1412];
   assign A[3][4][4]    = S_in[1476];
   assign A[4][4][4]    = S_in[1540];
   assign A[0][0][5]    = S_in[5];
   assign A[1][0][5]    = S_in[69];
   assign A[2][0][5]    = S_in[133];
   assign A[3][0][5]    = S_in[197];
   assign A[4][0][5]    = S_in[261];
   assign A[0][1][5]    = S_in[325];
   assign A[1][1][5]    = S_in[389];
   assign A[2][1][5]    = S_in[453];
   assign A[3][1][5]    = S_in[517];
   assign A[4][1][5]    = S_in[581];
   assign A[0][2][5]    = S_in[645];
   assign A[1][2][5]    = S_in[709];
   assign A[2][2][5]    = S_in[773];
   assign A[3][2][5]    = S_in[837];
   assign A[4][2][5]    = S_in[901];
   assign A[0][3][5]    = S_in[965];
   assign A[1][3][5]    = S_in[1029];
   assign A[2][3][5]    = S_in[1093];
   assign A[3][3][5]    = S_in[1157];
   assign A[4][3][5]    = S_in[1221];
   assign A[0][4][5]    = S_in[1285];
   assign A[1][4][5]    = S_in[1349];
   assign A[2][4][5]    = S_in[1413];
   assign A[3][4][5]    = S_in[1477];
   assign A[4][4][5]    = S_in[1541];
   assign A[0][0][6]    = S_in[6];
   assign A[1][0][6]    = S_in[70];
   assign A[2][0][6]    = S_in[134];
   assign A[3][0][6]    = S_in[198];
   assign A[4][0][6]    = S_in[262];
   assign A[0][1][6]    = S_in[326];
   assign A[1][1][6]    = S_in[390];
   assign A[2][1][6]    = S_in[454];
   assign A[3][1][6]    = S_in[518];
   assign A[4][1][6]    = S_in[582];
   assign A[0][2][6]    = S_in[646];
   assign A[1][2][6]    = S_in[710];
   assign A[2][2][6]    = S_in[774];
   assign A[3][2][6]    = S_in[838];
   assign A[4][2][6]    = S_in[902];
   assign A[0][3][6]    = S_in[966];
   assign A[1][3][6]    = S_in[1030];
   assign A[2][3][6]    = S_in[1094];
   assign A[3][3][6]    = S_in[1158];
   assign A[4][3][6]    = S_in[1222];
   assign A[0][4][6]    = S_in[1286];
   assign A[1][4][6]    = S_in[1350];
   assign A[2][4][6]    = S_in[1414];
   assign A[3][4][6]    = S_in[1478];
   assign A[4][4][6]    = S_in[1542];
   assign A[0][0][7]    = S_in[7];
   assign A[1][0][7]    = S_in[71];
   assign A[2][0][7]    = S_in[135];
   assign A[3][0][7]    = S_in[199];
   assign A[4][0][7]    = S_in[263];
   assign A[0][1][7]    = S_in[327];
   assign A[1][1][7]    = S_in[391];
   assign A[2][1][7]    = S_in[455];
   assign A[3][1][7]    = S_in[519];
   assign A[4][1][7]    = S_in[583];
   assign A[0][2][7]    = S_in[647];
   assign A[1][2][7]    = S_in[711];
   assign A[2][2][7]    = S_in[775];
   assign A[3][2][7]    = S_in[839];
   assign A[4][2][7]    = S_in[903];
   assign A[0][3][7]    = S_in[967];
   assign A[1][3][7]    = S_in[1031];
   assign A[2][3][7]    = S_in[1095];
   assign A[3][3][7]    = S_in[1159];
   assign A[4][3][7]    = S_in[1223];
   assign A[0][4][7]    = S_in[1287];
   assign A[1][4][7]    = S_in[1351];
   assign A[2][4][7]    = S_in[1415];
   assign A[3][4][7]    = S_in[1479];
   assign A[4][4][7]    = S_in[1543];
   assign A[0][0][8]    = S_in[8];
   assign A[1][0][8]    = S_in[72];
   assign A[2][0][8]    = S_in[136];
   assign A[3][0][8]    = S_in[200];
   assign A[4][0][8]    = S_in[264];
   assign A[0][1][8]    = S_in[328];
   assign A[1][1][8]    = S_in[392];
   assign A[2][1][8]    = S_in[456];
   assign A[3][1][8]    = S_in[520];
   assign A[4][1][8]    = S_in[584];
   assign A[0][2][8]    = S_in[648];
   assign A[1][2][8]    = S_in[712];
   assign A[2][2][8]    = S_in[776];
   assign A[3][2][8]    = S_in[840];
   assign A[4][2][8]    = S_in[904];
   assign A[0][3][8]    = S_in[968];
   assign A[1][3][8]    = S_in[1032];
   assign A[2][3][8]    = S_in[1096];
   assign A[3][3][8]    = S_in[1160];
   assign A[4][3][8]    = S_in[1224];
   assign A[0][4][8]    = S_in[1288];
   assign A[1][4][8]    = S_in[1352];
   assign A[2][4][8]    = S_in[1416];
   assign A[3][4][8]    = S_in[1480];
   assign A[4][4][8]    = S_in[1544];
   assign A[0][0][9]    = S_in[9];
   assign A[1][0][9]    = S_in[73];
   assign A[2][0][9]    = S_in[137];
   assign A[3][0][9]    = S_in[201];
   assign A[4][0][9]    = S_in[265];
   assign A[0][1][9]    = S_in[329];
   assign A[1][1][9]    = S_in[393];
   assign A[2][1][9]    = S_in[457];
   assign A[3][1][9]    = S_in[521];
   assign A[4][1][9]    = S_in[585];
   assign A[0][2][9]    = S_in[649];
   assign A[1][2][9]    = S_in[713];
   assign A[2][2][9]    = S_in[777];
   assign A[3][2][9]    = S_in[841];
   assign A[4][2][9]    = S_in[905];
   assign A[0][3][9]    = S_in[969];
   assign A[1][3][9]    = S_in[1033];
   assign A[2][3][9]    = S_in[1097];
   assign A[3][3][9]    = S_in[1161];
   assign A[4][3][9]    = S_in[1225];
   assign A[0][4][9]    = S_in[1289];
   assign A[1][4][9]    = S_in[1353];
   assign A[2][4][9]    = S_in[1417];
   assign A[3][4][9]    = S_in[1481];
   assign A[4][4][9]    = S_in[1545];
   assign A[0][0][10]    = S_in[10];
   assign A[1][0][10]    = S_in[74];
   assign A[2][0][10]    = S_in[138];
   assign A[3][0][10]    = S_in[202];
   assign A[4][0][10]    = S_in[266];
   assign A[0][1][10]    = S_in[330];
   assign A[1][1][10]    = S_in[394];
   assign A[2][1][10]    = S_in[458];
   assign A[3][1][10]    = S_in[522];
   assign A[4][1][10]    = S_in[586];
   assign A[0][2][10]    = S_in[650];
   assign A[1][2][10]    = S_in[714];
   assign A[2][2][10]    = S_in[778];
   assign A[3][2][10]    = S_in[842];
   assign A[4][2][10]    = S_in[906];
   assign A[0][3][10]    = S_in[970];
   assign A[1][3][10]    = S_in[1034];
   assign A[2][3][10]    = S_in[1098];
   assign A[3][3][10]    = S_in[1162];
   assign A[4][3][10]    = S_in[1226];
   assign A[0][4][10]    = S_in[1290];
   assign A[1][4][10]    = S_in[1354];
   assign A[2][4][10]    = S_in[1418];
   assign A[3][4][10]    = S_in[1482];
   assign A[4][4][10]    = S_in[1546];
   assign A[0][0][11]    = S_in[11];
   assign A[1][0][11]    = S_in[75];
   assign A[2][0][11]    = S_in[139];
   assign A[3][0][11]    = S_in[203];
   assign A[4][0][11]    = S_in[267];
   assign A[0][1][11]    = S_in[331];
   assign A[1][1][11]    = S_in[395];
   assign A[2][1][11]    = S_in[459];
   assign A[3][1][11]    = S_in[523];
   assign A[4][1][11]    = S_in[587];
   assign A[0][2][11]    = S_in[651];
   assign A[1][2][11]    = S_in[715];
   assign A[2][2][11]    = S_in[779];
   assign A[3][2][11]    = S_in[843];
   assign A[4][2][11]    = S_in[907];
   assign A[0][3][11]    = S_in[971];
   assign A[1][3][11]    = S_in[1035];
   assign A[2][3][11]    = S_in[1099];
   assign A[3][3][11]    = S_in[1163];
   assign A[4][3][11]    = S_in[1227];
   assign A[0][4][11]    = S_in[1291];
   assign A[1][4][11]    = S_in[1355];
   assign A[2][4][11]    = S_in[1419];
   assign A[3][4][11]    = S_in[1483];
   assign A[4][4][11]    = S_in[1547];
   assign A[0][0][12]    = S_in[12];
   assign A[1][0][12]    = S_in[76];
   assign A[2][0][12]    = S_in[140];
   assign A[3][0][12]    = S_in[204];
   assign A[4][0][12]    = S_in[268];
   assign A[0][1][12]    = S_in[332];
   assign A[1][1][12]    = S_in[396];
   assign A[2][1][12]    = S_in[460];
   assign A[3][1][12]    = S_in[524];
   assign A[4][1][12]    = S_in[588];
   assign A[0][2][12]    = S_in[652];
   assign A[1][2][12]    = S_in[716];
   assign A[2][2][12]    = S_in[780];
   assign A[3][2][12]    = S_in[844];
   assign A[4][2][12]    = S_in[908];
   assign A[0][3][12]    = S_in[972];
   assign A[1][3][12]    = S_in[1036];
   assign A[2][3][12]    = S_in[1100];
   assign A[3][3][12]    = S_in[1164];
   assign A[4][3][12]    = S_in[1228];
   assign A[0][4][12]    = S_in[1292];
   assign A[1][4][12]    = S_in[1356];
   assign A[2][4][12]    = S_in[1420];
   assign A[3][4][12]    = S_in[1484];
   assign A[4][4][12]    = S_in[1548];
   assign A[0][0][13]    = S_in[13];
   assign A[1][0][13]    = S_in[77];
   assign A[2][0][13]    = S_in[141];
   assign A[3][0][13]    = S_in[205];
   assign A[4][0][13]    = S_in[269];
   assign A[0][1][13]    = S_in[333];
   assign A[1][1][13]    = S_in[397];
   assign A[2][1][13]    = S_in[461];
   assign A[3][1][13]    = S_in[525];
   assign A[4][1][13]    = S_in[589];
   assign A[0][2][13]    = S_in[653];
   assign A[1][2][13]    = S_in[717];
   assign A[2][2][13]    = S_in[781];
   assign A[3][2][13]    = S_in[845];
   assign A[4][2][13]    = S_in[909];
   assign A[0][3][13]    = S_in[973];
   assign A[1][3][13]    = S_in[1037];
   assign A[2][3][13]    = S_in[1101];
   assign A[3][3][13]    = S_in[1165];
   assign A[4][3][13]    = S_in[1229];
   assign A[0][4][13]    = S_in[1293];
   assign A[1][4][13]    = S_in[1357];
   assign A[2][4][13]    = S_in[1421];
   assign A[3][4][13]    = S_in[1485];
   assign A[4][4][13]    = S_in[1549];
   assign A[0][0][14]    = S_in[14];
   assign A[1][0][14]    = S_in[78];
   assign A[2][0][14]    = S_in[142];
   assign A[3][0][14]    = S_in[206];
   assign A[4][0][14]    = S_in[270];
   assign A[0][1][14]    = S_in[334];
   assign A[1][1][14]    = S_in[398];
   assign A[2][1][14]    = S_in[462];
   assign A[3][1][14]    = S_in[526];
   assign A[4][1][14]    = S_in[590];
   assign A[0][2][14]    = S_in[654];
   assign A[1][2][14]    = S_in[718];
   assign A[2][2][14]    = S_in[782];
   assign A[3][2][14]    = S_in[846];
   assign A[4][2][14]    = S_in[910];
   assign A[0][3][14]    = S_in[974];
   assign A[1][3][14]    = S_in[1038];
   assign A[2][3][14]    = S_in[1102];
   assign A[3][3][14]    = S_in[1166];
   assign A[4][3][14]    = S_in[1230];
   assign A[0][4][14]    = S_in[1294];
   assign A[1][4][14]    = S_in[1358];
   assign A[2][4][14]    = S_in[1422];
   assign A[3][4][14]    = S_in[1486];
   assign A[4][4][14]    = S_in[1550];
   assign A[0][0][15]    = S_in[15];
   assign A[1][0][15]    = S_in[79];
   assign A[2][0][15]    = S_in[143];
   assign A[3][0][15]    = S_in[207];
   assign A[4][0][15]    = S_in[271];
   assign A[0][1][15]    = S_in[335];
   assign A[1][1][15]    = S_in[399];
   assign A[2][1][15]    = S_in[463];
   assign A[3][1][15]    = S_in[527];
   assign A[4][1][15]    = S_in[591];
   assign A[0][2][15]    = S_in[655];
   assign A[1][2][15]    = S_in[719];
   assign A[2][2][15]    = S_in[783];
   assign A[3][2][15]    = S_in[847];
   assign A[4][2][15]    = S_in[911];
   assign A[0][3][15]    = S_in[975];
   assign A[1][3][15]    = S_in[1039];
   assign A[2][3][15]    = S_in[1103];
   assign A[3][3][15]    = S_in[1167];
   assign A[4][3][15]    = S_in[1231];
   assign A[0][4][15]    = S_in[1295];
   assign A[1][4][15]    = S_in[1359];
   assign A[2][4][15]    = S_in[1423];
   assign A[3][4][15]    = S_in[1487];
   assign A[4][4][15]    = S_in[1551];
   assign A[0][0][16]    = S_in[16];
   assign A[1][0][16]    = S_in[80];
   assign A[2][0][16]    = S_in[144];
   assign A[3][0][16]    = S_in[208];
   assign A[4][0][16]    = S_in[272];
   assign A[0][1][16]    = S_in[336];
   assign A[1][1][16]    = S_in[400];
   assign A[2][1][16]    = S_in[464];
   assign A[3][1][16]    = S_in[528];
   assign A[4][1][16]    = S_in[592];
   assign A[0][2][16]    = S_in[656];
   assign A[1][2][16]    = S_in[720];
   assign A[2][2][16]    = S_in[784];
   assign A[3][2][16]    = S_in[848];
   assign A[4][2][16]    = S_in[912];
   assign A[0][3][16]    = S_in[976];
   assign A[1][3][16]    = S_in[1040];
   assign A[2][3][16]    = S_in[1104];
   assign A[3][3][16]    = S_in[1168];
   assign A[4][3][16]    = S_in[1232];
   assign A[0][4][16]    = S_in[1296];
   assign A[1][4][16]    = S_in[1360];
   assign A[2][4][16]    = S_in[1424];
   assign A[3][4][16]    = S_in[1488];
   assign A[4][4][16]    = S_in[1552];
   assign A[0][0][17]    = S_in[17];
   assign A[1][0][17]    = S_in[81];
   assign A[2][0][17]    = S_in[145];
   assign A[3][0][17]    = S_in[209];
   assign A[4][0][17]    = S_in[273];
   assign A[0][1][17]    = S_in[337];
   assign A[1][1][17]    = S_in[401];
   assign A[2][1][17]    = S_in[465];
   assign A[3][1][17]    = S_in[529];
   assign A[4][1][17]    = S_in[593];
   assign A[0][2][17]    = S_in[657];
   assign A[1][2][17]    = S_in[721];
   assign A[2][2][17]    = S_in[785];
   assign A[3][2][17]    = S_in[849];
   assign A[4][2][17]    = S_in[913];
   assign A[0][3][17]    = S_in[977];
   assign A[1][3][17]    = S_in[1041];
   assign A[2][3][17]    = S_in[1105];
   assign A[3][3][17]    = S_in[1169];
   assign A[4][3][17]    = S_in[1233];
   assign A[0][4][17]    = S_in[1297];
   assign A[1][4][17]    = S_in[1361];
   assign A[2][4][17]    = S_in[1425];
   assign A[3][4][17]    = S_in[1489];
   assign A[4][4][17]    = S_in[1553];
   assign A[0][0][18]    = S_in[18];
   assign A[1][0][18]    = S_in[82];
   assign A[2][0][18]    = S_in[146];
   assign A[3][0][18]    = S_in[210];
   assign A[4][0][18]    = S_in[274];
   assign A[0][1][18]    = S_in[338];
   assign A[1][1][18]    = S_in[402];
   assign A[2][1][18]    = S_in[466];
   assign A[3][1][18]    = S_in[530];
   assign A[4][1][18]    = S_in[594];
   assign A[0][2][18]    = S_in[658];
   assign A[1][2][18]    = S_in[722];
   assign A[2][2][18]    = S_in[786];
   assign A[3][2][18]    = S_in[850];
   assign A[4][2][18]    = S_in[914];
   assign A[0][3][18]    = S_in[978];
   assign A[1][3][18]    = S_in[1042];
   assign A[2][3][18]    = S_in[1106];
   assign A[3][3][18]    = S_in[1170];
   assign A[4][3][18]    = S_in[1234];
   assign A[0][4][18]    = S_in[1298];
   assign A[1][4][18]    = S_in[1362];
   assign A[2][4][18]    = S_in[1426];
   assign A[3][4][18]    = S_in[1490];
   assign A[4][4][18]    = S_in[1554];
   assign A[0][0][19]    = S_in[19];
   assign A[1][0][19]    = S_in[83];
   assign A[2][0][19]    = S_in[147];
   assign A[3][0][19]    = S_in[211];
   assign A[4][0][19]    = S_in[275];
   assign A[0][1][19]    = S_in[339];
   assign A[1][1][19]    = S_in[403];
   assign A[2][1][19]    = S_in[467];
   assign A[3][1][19]    = S_in[531];
   assign A[4][1][19]    = S_in[595];
   assign A[0][2][19]    = S_in[659];
   assign A[1][2][19]    = S_in[723];
   assign A[2][2][19]    = S_in[787];
   assign A[3][2][19]    = S_in[851];
   assign A[4][2][19]    = S_in[915];
   assign A[0][3][19]    = S_in[979];
   assign A[1][3][19]    = S_in[1043];
   assign A[2][3][19]    = S_in[1107];
   assign A[3][3][19]    = S_in[1171];
   assign A[4][3][19]    = S_in[1235];
   assign A[0][4][19]    = S_in[1299];
   assign A[1][4][19]    = S_in[1363];
   assign A[2][4][19]    = S_in[1427];
   assign A[3][4][19]    = S_in[1491];
   assign A[4][4][19]    = S_in[1555];
   assign A[0][0][20]    = S_in[20];
   assign A[1][0][20]    = S_in[84];
   assign A[2][0][20]    = S_in[148];
   assign A[3][0][20]    = S_in[212];
   assign A[4][0][20]    = S_in[276];
   assign A[0][1][20]    = S_in[340];
   assign A[1][1][20]    = S_in[404];
   assign A[2][1][20]    = S_in[468];
   assign A[3][1][20]    = S_in[532];
   assign A[4][1][20]    = S_in[596];
   assign A[0][2][20]    = S_in[660];
   assign A[1][2][20]    = S_in[724];
   assign A[2][2][20]    = S_in[788];
   assign A[3][2][20]    = S_in[852];
   assign A[4][2][20]    = S_in[916];
   assign A[0][3][20]    = S_in[980];
   assign A[1][3][20]    = S_in[1044];
   assign A[2][3][20]    = S_in[1108];
   assign A[3][3][20]    = S_in[1172];
   assign A[4][3][20]    = S_in[1236];
   assign A[0][4][20]    = S_in[1300];
   assign A[1][4][20]    = S_in[1364];
   assign A[2][4][20]    = S_in[1428];
   assign A[3][4][20]    = S_in[1492];
   assign A[4][4][20]    = S_in[1556];
   assign A[0][0][21]    = S_in[21];
   assign A[1][0][21]    = S_in[85];
   assign A[2][0][21]    = S_in[149];
   assign A[3][0][21]    = S_in[213];
   assign A[4][0][21]    = S_in[277];
   assign A[0][1][21]    = S_in[341];
   assign A[1][1][21]    = S_in[405];
   assign A[2][1][21]    = S_in[469];
   assign A[3][1][21]    = S_in[533];
   assign A[4][1][21]    = S_in[597];
   assign A[0][2][21]    = S_in[661];
   assign A[1][2][21]    = S_in[725];
   assign A[2][2][21]    = S_in[789];
   assign A[3][2][21]    = S_in[853];
   assign A[4][2][21]    = S_in[917];
   assign A[0][3][21]    = S_in[981];
   assign A[1][3][21]    = S_in[1045];
   assign A[2][3][21]    = S_in[1109];
   assign A[3][3][21]    = S_in[1173];
   assign A[4][3][21]    = S_in[1237];
   assign A[0][4][21]    = S_in[1301];
   assign A[1][4][21]    = S_in[1365];
   assign A[2][4][21]    = S_in[1429];
   assign A[3][4][21]    = S_in[1493];
   assign A[4][4][21]    = S_in[1557];
   assign A[0][0][22]    = S_in[22];
   assign A[1][0][22]    = S_in[86];
   assign A[2][0][22]    = S_in[150];
   assign A[3][0][22]    = S_in[214];
   assign A[4][0][22]    = S_in[278];
   assign A[0][1][22]    = S_in[342];
   assign A[1][1][22]    = S_in[406];
   assign A[2][1][22]    = S_in[470];
   assign A[3][1][22]    = S_in[534];
   assign A[4][1][22]    = S_in[598];
   assign A[0][2][22]    = S_in[662];
   assign A[1][2][22]    = S_in[726];
   assign A[2][2][22]    = S_in[790];
   assign A[3][2][22]    = S_in[854];
   assign A[4][2][22]    = S_in[918];
   assign A[0][3][22]    = S_in[982];
   assign A[1][3][22]    = S_in[1046];
   assign A[2][3][22]    = S_in[1110];
   assign A[3][3][22]    = S_in[1174];
   assign A[4][3][22]    = S_in[1238];
   assign A[0][4][22]    = S_in[1302];
   assign A[1][4][22]    = S_in[1366];
   assign A[2][4][22]    = S_in[1430];
   assign A[3][4][22]    = S_in[1494];
   assign A[4][4][22]    = S_in[1558];
   assign A[0][0][23]    = S_in[23];
   assign A[1][0][23]    = S_in[87];
   assign A[2][0][23]    = S_in[151];
   assign A[3][0][23]    = S_in[215];
   assign A[4][0][23]    = S_in[279];
   assign A[0][1][23]    = S_in[343];
   assign A[1][1][23]    = S_in[407];
   assign A[2][1][23]    = S_in[471];
   assign A[3][1][23]    = S_in[535];
   assign A[4][1][23]    = S_in[599];
   assign A[0][2][23]    = S_in[663];
   assign A[1][2][23]    = S_in[727];
   assign A[2][2][23]    = S_in[791];
   assign A[3][2][23]    = S_in[855];
   assign A[4][2][23]    = S_in[919];
   assign A[0][3][23]    = S_in[983];
   assign A[1][3][23]    = S_in[1047];
   assign A[2][3][23]    = S_in[1111];
   assign A[3][3][23]    = S_in[1175];
   assign A[4][3][23]    = S_in[1239];
   assign A[0][4][23]    = S_in[1303];
   assign A[1][4][23]    = S_in[1367];
   assign A[2][4][23]    = S_in[1431];
   assign A[3][4][23]    = S_in[1495];
   assign A[4][4][23]    = S_in[1559];
   assign A[0][0][24]    = S_in[24];
   assign A[1][0][24]    = S_in[88];
   assign A[2][0][24]    = S_in[152];
   assign A[3][0][24]    = S_in[216];
   assign A[4][0][24]    = S_in[280];
   assign A[0][1][24]    = S_in[344];
   assign A[1][1][24]    = S_in[408];
   assign A[2][1][24]    = S_in[472];
   assign A[3][1][24]    = S_in[536];
   assign A[4][1][24]    = S_in[600];
   assign A[0][2][24]    = S_in[664];
   assign A[1][2][24]    = S_in[728];
   assign A[2][2][24]    = S_in[792];
   assign A[3][2][24]    = S_in[856];
   assign A[4][2][24]    = S_in[920];
   assign A[0][3][24]    = S_in[984];
   assign A[1][3][24]    = S_in[1048];
   assign A[2][3][24]    = S_in[1112];
   assign A[3][3][24]    = S_in[1176];
   assign A[4][3][24]    = S_in[1240];
   assign A[0][4][24]    = S_in[1304];
   assign A[1][4][24]    = S_in[1368];
   assign A[2][4][24]    = S_in[1432];
   assign A[3][4][24]    = S_in[1496];
   assign A[4][4][24]    = S_in[1560];
   assign A[0][0][25]    = S_in[25];
   assign A[1][0][25]    = S_in[89];
   assign A[2][0][25]    = S_in[153];
   assign A[3][0][25]    = S_in[217];
   assign A[4][0][25]    = S_in[281];
   assign A[0][1][25]    = S_in[345];
   assign A[1][1][25]    = S_in[409];
   assign A[2][1][25]    = S_in[473];
   assign A[3][1][25]    = S_in[537];
   assign A[4][1][25]    = S_in[601];
   assign A[0][2][25]    = S_in[665];
   assign A[1][2][25]    = S_in[729];
   assign A[2][2][25]    = S_in[793];
   assign A[3][2][25]    = S_in[857];
   assign A[4][2][25]    = S_in[921];
   assign A[0][3][25]    = S_in[985];
   assign A[1][3][25]    = S_in[1049];
   assign A[2][3][25]    = S_in[1113];
   assign A[3][3][25]    = S_in[1177];
   assign A[4][3][25]    = S_in[1241];
   assign A[0][4][25]    = S_in[1305];
   assign A[1][4][25]    = S_in[1369];
   assign A[2][4][25]    = S_in[1433];
   assign A[3][4][25]    = S_in[1497];
   assign A[4][4][25]    = S_in[1561];
   assign A[0][0][26]    = S_in[26];
   assign A[1][0][26]    = S_in[90];
   assign A[2][0][26]    = S_in[154];
   assign A[3][0][26]    = S_in[218];
   assign A[4][0][26]    = S_in[282];
   assign A[0][1][26]    = S_in[346];
   assign A[1][1][26]    = S_in[410];
   assign A[2][1][26]    = S_in[474];
   assign A[3][1][26]    = S_in[538];
   assign A[4][1][26]    = S_in[602];
   assign A[0][2][26]    = S_in[666];
   assign A[1][2][26]    = S_in[730];
   assign A[2][2][26]    = S_in[794];
   assign A[3][2][26]    = S_in[858];
   assign A[4][2][26]    = S_in[922];
   assign A[0][3][26]    = S_in[986];
   assign A[1][3][26]    = S_in[1050];
   assign A[2][3][26]    = S_in[1114];
   assign A[3][3][26]    = S_in[1178];
   assign A[4][3][26]    = S_in[1242];
   assign A[0][4][26]    = S_in[1306];
   assign A[1][4][26]    = S_in[1370];
   assign A[2][4][26]    = S_in[1434];
   assign A[3][4][26]    = S_in[1498];
   assign A[4][4][26]    = S_in[1562];
   assign A[0][0][27]    = S_in[27];
   assign A[1][0][27]    = S_in[91];
   assign A[2][0][27]    = S_in[155];
   assign A[3][0][27]    = S_in[219];
   assign A[4][0][27]    = S_in[283];
   assign A[0][1][27]    = S_in[347];
   assign A[1][1][27]    = S_in[411];
   assign A[2][1][27]    = S_in[475];
   assign A[3][1][27]    = S_in[539];
   assign A[4][1][27]    = S_in[603];
   assign A[0][2][27]    = S_in[667];
   assign A[1][2][27]    = S_in[731];
   assign A[2][2][27]    = S_in[795];
   assign A[3][2][27]    = S_in[859];
   assign A[4][2][27]    = S_in[923];
   assign A[0][3][27]    = S_in[987];
   assign A[1][3][27]    = S_in[1051];
   assign A[2][3][27]    = S_in[1115];
   assign A[3][3][27]    = S_in[1179];
   assign A[4][3][27]    = S_in[1243];
   assign A[0][4][27]    = S_in[1307];
   assign A[1][4][27]    = S_in[1371];
   assign A[2][4][27]    = S_in[1435];
   assign A[3][4][27]    = S_in[1499];
   assign A[4][4][27]    = S_in[1563];
   assign A[0][0][28]    = S_in[28];
   assign A[1][0][28]    = S_in[92];
   assign A[2][0][28]    = S_in[156];
   assign A[3][0][28]    = S_in[220];
   assign A[4][0][28]    = S_in[284];
   assign A[0][1][28]    = S_in[348];
   assign A[1][1][28]    = S_in[412];
   assign A[2][1][28]    = S_in[476];
   assign A[3][1][28]    = S_in[540];
   assign A[4][1][28]    = S_in[604];
   assign A[0][2][28]    = S_in[668];
   assign A[1][2][28]    = S_in[732];
   assign A[2][2][28]    = S_in[796];
   assign A[3][2][28]    = S_in[860];
   assign A[4][2][28]    = S_in[924];
   assign A[0][3][28]    = S_in[988];
   assign A[1][3][28]    = S_in[1052];
   assign A[2][3][28]    = S_in[1116];
   assign A[3][3][28]    = S_in[1180];
   assign A[4][3][28]    = S_in[1244];
   assign A[0][4][28]    = S_in[1308];
   assign A[1][4][28]    = S_in[1372];
   assign A[2][4][28]    = S_in[1436];
   assign A[3][4][28]    = S_in[1500];
   assign A[4][4][28]    = S_in[1564];
   assign A[0][0][29]    = S_in[29];
   assign A[1][0][29]    = S_in[93];
   assign A[2][0][29]    = S_in[157];
   assign A[3][0][29]    = S_in[221];
   assign A[4][0][29]    = S_in[285];
   assign A[0][1][29]    = S_in[349];
   assign A[1][1][29]    = S_in[413];
   assign A[2][1][29]    = S_in[477];
   assign A[3][1][29]    = S_in[541];
   assign A[4][1][29]    = S_in[605];
   assign A[0][2][29]    = S_in[669];
   assign A[1][2][29]    = S_in[733];
   assign A[2][2][29]    = S_in[797];
   assign A[3][2][29]    = S_in[861];
   assign A[4][2][29]    = S_in[925];
   assign A[0][3][29]    = S_in[989];
   assign A[1][3][29]    = S_in[1053];
   assign A[2][3][29]    = S_in[1117];
   assign A[3][3][29]    = S_in[1181];
   assign A[4][3][29]    = S_in[1245];
   assign A[0][4][29]    = S_in[1309];
   assign A[1][4][29]    = S_in[1373];
   assign A[2][4][29]    = S_in[1437];
   assign A[3][4][29]    = S_in[1501];
   assign A[4][4][29]    = S_in[1565];
   assign A[0][0][30]    = S_in[30];
   assign A[1][0][30]    = S_in[94];
   assign A[2][0][30]    = S_in[158];
   assign A[3][0][30]    = S_in[222];
   assign A[4][0][30]    = S_in[286];
   assign A[0][1][30]    = S_in[350];
   assign A[1][1][30]    = S_in[414];
   assign A[2][1][30]    = S_in[478];
   assign A[3][1][30]    = S_in[542];
   assign A[4][1][30]    = S_in[606];
   assign A[0][2][30]    = S_in[670];
   assign A[1][2][30]    = S_in[734];
   assign A[2][2][30]    = S_in[798];
   assign A[3][2][30]    = S_in[862];
   assign A[4][2][30]    = S_in[926];
   assign A[0][3][30]    = S_in[990];
   assign A[1][3][30]    = S_in[1054];
   assign A[2][3][30]    = S_in[1118];
   assign A[3][3][30]    = S_in[1182];
   assign A[4][3][30]    = S_in[1246];
   assign A[0][4][30]    = S_in[1310];
   assign A[1][4][30]    = S_in[1374];
   assign A[2][4][30]    = S_in[1438];
   assign A[3][4][30]    = S_in[1502];
   assign A[4][4][30]    = S_in[1566];
   assign A[0][0][31]    = S_in[31];
   assign A[1][0][31]    = S_in[95];
   assign A[2][0][31]    = S_in[159];
   assign A[3][0][31]    = S_in[223];
   assign A[4][0][31]    = S_in[287];
   assign A[0][1][31]    = S_in[351];
   assign A[1][1][31]    = S_in[415];
   assign A[2][1][31]    = S_in[479];
   assign A[3][1][31]    = S_in[543];
   assign A[4][1][31]    = S_in[607];
   assign A[0][2][31]    = S_in[671];
   assign A[1][2][31]    = S_in[735];
   assign A[2][2][31]    = S_in[799];
   assign A[3][2][31]    = S_in[863];
   assign A[4][2][31]    = S_in[927];
   assign A[0][3][31]    = S_in[991];
   assign A[1][3][31]    = S_in[1055];
   assign A[2][3][31]    = S_in[1119];
   assign A[3][3][31]    = S_in[1183];
   assign A[4][3][31]    = S_in[1247];
   assign A[0][4][31]    = S_in[1311];
   assign A[1][4][31]    = S_in[1375];
   assign A[2][4][31]    = S_in[1439];
   assign A[3][4][31]    = S_in[1503];
   assign A[4][4][31]    = S_in[1567];
   assign A[0][0][32]    = S_in[32];
   assign A[1][0][32]    = S_in[96];
   assign A[2][0][32]    = S_in[160];
   assign A[3][0][32]    = S_in[224];
   assign A[4][0][32]    = S_in[288];
   assign A[0][1][32]    = S_in[352];
   assign A[1][1][32]    = S_in[416];
   assign A[2][1][32]    = S_in[480];
   assign A[3][1][32]    = S_in[544];
   assign A[4][1][32]    = S_in[608];
   assign A[0][2][32]    = S_in[672];
   assign A[1][2][32]    = S_in[736];
   assign A[2][2][32]    = S_in[800];
   assign A[3][2][32]    = S_in[864];
   assign A[4][2][32]    = S_in[928];
   assign A[0][3][32]    = S_in[992];
   assign A[1][3][32]    = S_in[1056];
   assign A[2][3][32]    = S_in[1120];
   assign A[3][3][32]    = S_in[1184];
   assign A[4][3][32]    = S_in[1248];
   assign A[0][4][32]    = S_in[1312];
   assign A[1][4][32]    = S_in[1376];
   assign A[2][4][32]    = S_in[1440];
   assign A[3][4][32]    = S_in[1504];
   assign A[4][4][32]    = S_in[1568];
   assign A[0][0][33]    = S_in[33];
   assign A[1][0][33]    = S_in[97];
   assign A[2][0][33]    = S_in[161];
   assign A[3][0][33]    = S_in[225];
   assign A[4][0][33]    = S_in[289];
   assign A[0][1][33]    = S_in[353];
   assign A[1][1][33]    = S_in[417];
   assign A[2][1][33]    = S_in[481];
   assign A[3][1][33]    = S_in[545];
   assign A[4][1][33]    = S_in[609];
   assign A[0][2][33]    = S_in[673];
   assign A[1][2][33]    = S_in[737];
   assign A[2][2][33]    = S_in[801];
   assign A[3][2][33]    = S_in[865];
   assign A[4][2][33]    = S_in[929];
   assign A[0][3][33]    = S_in[993];
   assign A[1][3][33]    = S_in[1057];
   assign A[2][3][33]    = S_in[1121];
   assign A[3][3][33]    = S_in[1185];
   assign A[4][3][33]    = S_in[1249];
   assign A[0][4][33]    = S_in[1313];
   assign A[1][4][33]    = S_in[1377];
   assign A[2][4][33]    = S_in[1441];
   assign A[3][4][33]    = S_in[1505];
   assign A[4][4][33]    = S_in[1569];
   assign A[0][0][34]    = S_in[34];
   assign A[1][0][34]    = S_in[98];
   assign A[2][0][34]    = S_in[162];
   assign A[3][0][34]    = S_in[226];
   assign A[4][0][34]    = S_in[290];
   assign A[0][1][34]    = S_in[354];
   assign A[1][1][34]    = S_in[418];
   assign A[2][1][34]    = S_in[482];
   assign A[3][1][34]    = S_in[546];
   assign A[4][1][34]    = S_in[610];
   assign A[0][2][34]    = S_in[674];
   assign A[1][2][34]    = S_in[738];
   assign A[2][2][34]    = S_in[802];
   assign A[3][2][34]    = S_in[866];
   assign A[4][2][34]    = S_in[930];
   assign A[0][3][34]    = S_in[994];
   assign A[1][3][34]    = S_in[1058];
   assign A[2][3][34]    = S_in[1122];
   assign A[3][3][34]    = S_in[1186];
   assign A[4][3][34]    = S_in[1250];
   assign A[0][4][34]    = S_in[1314];
   assign A[1][4][34]    = S_in[1378];
   assign A[2][4][34]    = S_in[1442];
   assign A[3][4][34]    = S_in[1506];
   assign A[4][4][34]    = S_in[1570];
   assign A[0][0][35]    = S_in[35];
   assign A[1][0][35]    = S_in[99];
   assign A[2][0][35]    = S_in[163];
   assign A[3][0][35]    = S_in[227];
   assign A[4][0][35]    = S_in[291];
   assign A[0][1][35]    = S_in[355];
   assign A[1][1][35]    = S_in[419];
   assign A[2][1][35]    = S_in[483];
   assign A[3][1][35]    = S_in[547];
   assign A[4][1][35]    = S_in[611];
   assign A[0][2][35]    = S_in[675];
   assign A[1][2][35]    = S_in[739];
   assign A[2][2][35]    = S_in[803];
   assign A[3][2][35]    = S_in[867];
   assign A[4][2][35]    = S_in[931];
   assign A[0][3][35]    = S_in[995];
   assign A[1][3][35]    = S_in[1059];
   assign A[2][3][35]    = S_in[1123];
   assign A[3][3][35]    = S_in[1187];
   assign A[4][3][35]    = S_in[1251];
   assign A[0][4][35]    = S_in[1315];
   assign A[1][4][35]    = S_in[1379];
   assign A[2][4][35]    = S_in[1443];
   assign A[3][4][35]    = S_in[1507];
   assign A[4][4][35]    = S_in[1571];
   assign A[0][0][36]    = S_in[36];
   assign A[1][0][36]    = S_in[100];
   assign A[2][0][36]    = S_in[164];
   assign A[3][0][36]    = S_in[228];
   assign A[4][0][36]    = S_in[292];
   assign A[0][1][36]    = S_in[356];
   assign A[1][1][36]    = S_in[420];
   assign A[2][1][36]    = S_in[484];
   assign A[3][1][36]    = S_in[548];
   assign A[4][1][36]    = S_in[612];
   assign A[0][2][36]    = S_in[676];
   assign A[1][2][36]    = S_in[740];
   assign A[2][2][36]    = S_in[804];
   assign A[3][2][36]    = S_in[868];
   assign A[4][2][36]    = S_in[932];
   assign A[0][3][36]    = S_in[996];
   assign A[1][3][36]    = S_in[1060];
   assign A[2][3][36]    = S_in[1124];
   assign A[3][3][36]    = S_in[1188];
   assign A[4][3][36]    = S_in[1252];
   assign A[0][4][36]    = S_in[1316];
   assign A[1][4][36]    = S_in[1380];
   assign A[2][4][36]    = S_in[1444];
   assign A[3][4][36]    = S_in[1508];
   assign A[4][4][36]    = S_in[1572];
   assign A[0][0][37]    = S_in[37];
   assign A[1][0][37]    = S_in[101];
   assign A[2][0][37]    = S_in[165];
   assign A[3][0][37]    = S_in[229];
   assign A[4][0][37]    = S_in[293];
   assign A[0][1][37]    = S_in[357];
   assign A[1][1][37]    = S_in[421];
   assign A[2][1][37]    = S_in[485];
   assign A[3][1][37]    = S_in[549];
   assign A[4][1][37]    = S_in[613];
   assign A[0][2][37]    = S_in[677];
   assign A[1][2][37]    = S_in[741];
   assign A[2][2][37]    = S_in[805];
   assign A[3][2][37]    = S_in[869];
   assign A[4][2][37]    = S_in[933];
   assign A[0][3][37]    = S_in[997];
   assign A[1][3][37]    = S_in[1061];
   assign A[2][3][37]    = S_in[1125];
   assign A[3][3][37]    = S_in[1189];
   assign A[4][3][37]    = S_in[1253];
   assign A[0][4][37]    = S_in[1317];
   assign A[1][4][37]    = S_in[1381];
   assign A[2][4][37]    = S_in[1445];
   assign A[3][4][37]    = S_in[1509];
   assign A[4][4][37]    = S_in[1573];
   assign A[0][0][38]    = S_in[38];
   assign A[1][0][38]    = S_in[102];
   assign A[2][0][38]    = S_in[166];
   assign A[3][0][38]    = S_in[230];
   assign A[4][0][38]    = S_in[294];
   assign A[0][1][38]    = S_in[358];
   assign A[1][1][38]    = S_in[422];
   assign A[2][1][38]    = S_in[486];
   assign A[3][1][38]    = S_in[550];
   assign A[4][1][38]    = S_in[614];
   assign A[0][2][38]    = S_in[678];
   assign A[1][2][38]    = S_in[742];
   assign A[2][2][38]    = S_in[806];
   assign A[3][2][38]    = S_in[870];
   assign A[4][2][38]    = S_in[934];
   assign A[0][3][38]    = S_in[998];
   assign A[1][3][38]    = S_in[1062];
   assign A[2][3][38]    = S_in[1126];
   assign A[3][3][38]    = S_in[1190];
   assign A[4][3][38]    = S_in[1254];
   assign A[0][4][38]    = S_in[1318];
   assign A[1][4][38]    = S_in[1382];
   assign A[2][4][38]    = S_in[1446];
   assign A[3][4][38]    = S_in[1510];
   assign A[4][4][38]    = S_in[1574];
   assign A[0][0][39]    = S_in[39];
   assign A[1][0][39]    = S_in[103];
   assign A[2][0][39]    = S_in[167];
   assign A[3][0][39]    = S_in[231];
   assign A[4][0][39]    = S_in[295];
   assign A[0][1][39]    = S_in[359];
   assign A[1][1][39]    = S_in[423];
   assign A[2][1][39]    = S_in[487];
   assign A[3][1][39]    = S_in[551];
   assign A[4][1][39]    = S_in[615];
   assign A[0][2][39]    = S_in[679];
   assign A[1][2][39]    = S_in[743];
   assign A[2][2][39]    = S_in[807];
   assign A[3][2][39]    = S_in[871];
   assign A[4][2][39]    = S_in[935];
   assign A[0][3][39]    = S_in[999];
   assign A[1][3][39]    = S_in[1063];
   assign A[2][3][39]    = S_in[1127];
   assign A[3][3][39]    = S_in[1191];
   assign A[4][3][39]    = S_in[1255];
   assign A[0][4][39]    = S_in[1319];
   assign A[1][4][39]    = S_in[1383];
   assign A[2][4][39]    = S_in[1447];
   assign A[3][4][39]    = S_in[1511];
   assign A[4][4][39]    = S_in[1575];
   assign A[0][0][40]    = S_in[40];
   assign A[1][0][40]    = S_in[104];
   assign A[2][0][40]    = S_in[168];
   assign A[3][0][40]    = S_in[232];
   assign A[4][0][40]    = S_in[296];
   assign A[0][1][40]    = S_in[360];
   assign A[1][1][40]    = S_in[424];
   assign A[2][1][40]    = S_in[488];
   assign A[3][1][40]    = S_in[552];
   assign A[4][1][40]    = S_in[616];
   assign A[0][2][40]    = S_in[680];
   assign A[1][2][40]    = S_in[744];
   assign A[2][2][40]    = S_in[808];
   assign A[3][2][40]    = S_in[872];
   assign A[4][2][40]    = S_in[936];
   assign A[0][3][40]    = S_in[1000];
   assign A[1][3][40]    = S_in[1064];
   assign A[2][3][40]    = S_in[1128];
   assign A[3][3][40]    = S_in[1192];
   assign A[4][3][40]    = S_in[1256];
   assign A[0][4][40]    = S_in[1320];
   assign A[1][4][40]    = S_in[1384];
   assign A[2][4][40]    = S_in[1448];
   assign A[3][4][40]    = S_in[1512];
   assign A[4][4][40]    = S_in[1576];
   assign A[0][0][41]    = S_in[41];
   assign A[1][0][41]    = S_in[105];
   assign A[2][0][41]    = S_in[169];
   assign A[3][0][41]    = S_in[233];
   assign A[4][0][41]    = S_in[297];
   assign A[0][1][41]    = S_in[361];
   assign A[1][1][41]    = S_in[425];
   assign A[2][1][41]    = S_in[489];
   assign A[3][1][41]    = S_in[553];
   assign A[4][1][41]    = S_in[617];
   assign A[0][2][41]    = S_in[681];
   assign A[1][2][41]    = S_in[745];
   assign A[2][2][41]    = S_in[809];
   assign A[3][2][41]    = S_in[873];
   assign A[4][2][41]    = S_in[937];
   assign A[0][3][41]    = S_in[1001];
   assign A[1][3][41]    = S_in[1065];
   assign A[2][3][41]    = S_in[1129];
   assign A[3][3][41]    = S_in[1193];
   assign A[4][3][41]    = S_in[1257];
   assign A[0][4][41]    = S_in[1321];
   assign A[1][4][41]    = S_in[1385];
   assign A[2][4][41]    = S_in[1449];
   assign A[3][4][41]    = S_in[1513];
   assign A[4][4][41]    = S_in[1577];
   assign A[0][0][42]    = S_in[42];
   assign A[1][0][42]    = S_in[106];
   assign A[2][0][42]    = S_in[170];
   assign A[3][0][42]    = S_in[234];
   assign A[4][0][42]    = S_in[298];
   assign A[0][1][42]    = S_in[362];
   assign A[1][1][42]    = S_in[426];
   assign A[2][1][42]    = S_in[490];
   assign A[3][1][42]    = S_in[554];
   assign A[4][1][42]    = S_in[618];
   assign A[0][2][42]    = S_in[682];
   assign A[1][2][42]    = S_in[746];
   assign A[2][2][42]    = S_in[810];
   assign A[3][2][42]    = S_in[874];
   assign A[4][2][42]    = S_in[938];
   assign A[0][3][42]    = S_in[1002];
   assign A[1][3][42]    = S_in[1066];
   assign A[2][3][42]    = S_in[1130];
   assign A[3][3][42]    = S_in[1194];
   assign A[4][3][42]    = S_in[1258];
   assign A[0][4][42]    = S_in[1322];
   assign A[1][4][42]    = S_in[1386];
   assign A[2][4][42]    = S_in[1450];
   assign A[3][4][42]    = S_in[1514];
   assign A[4][4][42]    = S_in[1578];
   assign A[0][0][43]    = S_in[43];
   assign A[1][0][43]    = S_in[107];
   assign A[2][0][43]    = S_in[171];
   assign A[3][0][43]    = S_in[235];
   assign A[4][0][43]    = S_in[299];
   assign A[0][1][43]    = S_in[363];
   assign A[1][1][43]    = S_in[427];
   assign A[2][1][43]    = S_in[491];
   assign A[3][1][43]    = S_in[555];
   assign A[4][1][43]    = S_in[619];
   assign A[0][2][43]    = S_in[683];
   assign A[1][2][43]    = S_in[747];
   assign A[2][2][43]    = S_in[811];
   assign A[3][2][43]    = S_in[875];
   assign A[4][2][43]    = S_in[939];
   assign A[0][3][43]    = S_in[1003];
   assign A[1][3][43]    = S_in[1067];
   assign A[2][3][43]    = S_in[1131];
   assign A[3][3][43]    = S_in[1195];
   assign A[4][3][43]    = S_in[1259];
   assign A[0][4][43]    = S_in[1323];
   assign A[1][4][43]    = S_in[1387];
   assign A[2][4][43]    = S_in[1451];
   assign A[3][4][43]    = S_in[1515];
   assign A[4][4][43]    = S_in[1579];
   assign A[0][0][44]    = S_in[44];
   assign A[1][0][44]    = S_in[108];
   assign A[2][0][44]    = S_in[172];
   assign A[3][0][44]    = S_in[236];
   assign A[4][0][44]    = S_in[300];
   assign A[0][1][44]    = S_in[364];
   assign A[1][1][44]    = S_in[428];
   assign A[2][1][44]    = S_in[492];
   assign A[3][1][44]    = S_in[556];
   assign A[4][1][44]    = S_in[620];
   assign A[0][2][44]    = S_in[684];
   assign A[1][2][44]    = S_in[748];
   assign A[2][2][44]    = S_in[812];
   assign A[3][2][44]    = S_in[876];
   assign A[4][2][44]    = S_in[940];
   assign A[0][3][44]    = S_in[1004];
   assign A[1][3][44]    = S_in[1068];
   assign A[2][3][44]    = S_in[1132];
   assign A[3][3][44]    = S_in[1196];
   assign A[4][3][44]    = S_in[1260];
   assign A[0][4][44]    = S_in[1324];
   assign A[1][4][44]    = S_in[1388];
   assign A[2][4][44]    = S_in[1452];
   assign A[3][4][44]    = S_in[1516];
   assign A[4][4][44]    = S_in[1580];
   assign A[0][0][45]    = S_in[45];
   assign A[1][0][45]    = S_in[109];
   assign A[2][0][45]    = S_in[173];
   assign A[3][0][45]    = S_in[237];
   assign A[4][0][45]    = S_in[301];
   assign A[0][1][45]    = S_in[365];
   assign A[1][1][45]    = S_in[429];
   assign A[2][1][45]    = S_in[493];
   assign A[3][1][45]    = S_in[557];
   assign A[4][1][45]    = S_in[621];
   assign A[0][2][45]    = S_in[685];
   assign A[1][2][45]    = S_in[749];
   assign A[2][2][45]    = S_in[813];
   assign A[3][2][45]    = S_in[877];
   assign A[4][2][45]    = S_in[941];
   assign A[0][3][45]    = S_in[1005];
   assign A[1][3][45]    = S_in[1069];
   assign A[2][3][45]    = S_in[1133];
   assign A[3][3][45]    = S_in[1197];
   assign A[4][3][45]    = S_in[1261];
   assign A[0][4][45]    = S_in[1325];
   assign A[1][4][45]    = S_in[1389];
   assign A[2][4][45]    = S_in[1453];
   assign A[3][4][45]    = S_in[1517];
   assign A[4][4][45]    = S_in[1581];
   assign A[0][0][46]    = S_in[46];
   assign A[1][0][46]    = S_in[110];
   assign A[2][0][46]    = S_in[174];
   assign A[3][0][46]    = S_in[238];
   assign A[4][0][46]    = S_in[302];
   assign A[0][1][46]    = S_in[366];
   assign A[1][1][46]    = S_in[430];
   assign A[2][1][46]    = S_in[494];
   assign A[3][1][46]    = S_in[558];
   assign A[4][1][46]    = S_in[622];
   assign A[0][2][46]    = S_in[686];
   assign A[1][2][46]    = S_in[750];
   assign A[2][2][46]    = S_in[814];
   assign A[3][2][46]    = S_in[878];
   assign A[4][2][46]    = S_in[942];
   assign A[0][3][46]    = S_in[1006];
   assign A[1][3][46]    = S_in[1070];
   assign A[2][3][46]    = S_in[1134];
   assign A[3][3][46]    = S_in[1198];
   assign A[4][3][46]    = S_in[1262];
   assign A[0][4][46]    = S_in[1326];
   assign A[1][4][46]    = S_in[1390];
   assign A[2][4][46]    = S_in[1454];
   assign A[3][4][46]    = S_in[1518];
   assign A[4][4][46]    = S_in[1582];
   assign A[0][0][47]    = S_in[47];
   assign A[1][0][47]    = S_in[111];
   assign A[2][0][47]    = S_in[175];
   assign A[3][0][47]    = S_in[239];
   assign A[4][0][47]    = S_in[303];
   assign A[0][1][47]    = S_in[367];
   assign A[1][1][47]    = S_in[431];
   assign A[2][1][47]    = S_in[495];
   assign A[3][1][47]    = S_in[559];
   assign A[4][1][47]    = S_in[623];
   assign A[0][2][47]    = S_in[687];
   assign A[1][2][47]    = S_in[751];
   assign A[2][2][47]    = S_in[815];
   assign A[3][2][47]    = S_in[879];
   assign A[4][2][47]    = S_in[943];
   assign A[0][3][47]    = S_in[1007];
   assign A[1][3][47]    = S_in[1071];
   assign A[2][3][47]    = S_in[1135];
   assign A[3][3][47]    = S_in[1199];
   assign A[4][3][47]    = S_in[1263];
   assign A[0][4][47]    = S_in[1327];
   assign A[1][4][47]    = S_in[1391];
   assign A[2][4][47]    = S_in[1455];
   assign A[3][4][47]    = S_in[1519];
   assign A[4][4][47]    = S_in[1583];
   assign A[0][0][48]    = S_in[48];
   assign A[1][0][48]    = S_in[112];
   assign A[2][0][48]    = S_in[176];
   assign A[3][0][48]    = S_in[240];
   assign A[4][0][48]    = S_in[304];
   assign A[0][1][48]    = S_in[368];
   assign A[1][1][48]    = S_in[432];
   assign A[2][1][48]    = S_in[496];
   assign A[3][1][48]    = S_in[560];
   assign A[4][1][48]    = S_in[624];
   assign A[0][2][48]    = S_in[688];
   assign A[1][2][48]    = S_in[752];
   assign A[2][2][48]    = S_in[816];
   assign A[3][2][48]    = S_in[880];
   assign A[4][2][48]    = S_in[944];
   assign A[0][3][48]    = S_in[1008];
   assign A[1][3][48]    = S_in[1072];
   assign A[2][3][48]    = S_in[1136];
   assign A[3][3][48]    = S_in[1200];
   assign A[4][3][48]    = S_in[1264];
   assign A[0][4][48]    = S_in[1328];
   assign A[1][4][48]    = S_in[1392];
   assign A[2][4][48]    = S_in[1456];
   assign A[3][4][48]    = S_in[1520];
   assign A[4][4][48]    = S_in[1584];
   assign A[0][0][49]    = S_in[49];
   assign A[1][0][49]    = S_in[113];
   assign A[2][0][49]    = S_in[177];
   assign A[3][0][49]    = S_in[241];
   assign A[4][0][49]    = S_in[305];
   assign A[0][1][49]    = S_in[369];
   assign A[1][1][49]    = S_in[433];
   assign A[2][1][49]    = S_in[497];
   assign A[3][1][49]    = S_in[561];
   assign A[4][1][49]    = S_in[625];
   assign A[0][2][49]    = S_in[689];
   assign A[1][2][49]    = S_in[753];
   assign A[2][2][49]    = S_in[817];
   assign A[3][2][49]    = S_in[881];
   assign A[4][2][49]    = S_in[945];
   assign A[0][3][49]    = S_in[1009];
   assign A[1][3][49]    = S_in[1073];
   assign A[2][3][49]    = S_in[1137];
   assign A[3][3][49]    = S_in[1201];
   assign A[4][3][49]    = S_in[1265];
   assign A[0][4][49]    = S_in[1329];
   assign A[1][4][49]    = S_in[1393];
   assign A[2][4][49]    = S_in[1457];
   assign A[3][4][49]    = S_in[1521];
   assign A[4][4][49]    = S_in[1585];
   assign A[0][0][50]    = S_in[50];
   assign A[1][0][50]    = S_in[114];
   assign A[2][0][50]    = S_in[178];
   assign A[3][0][50]    = S_in[242];
   assign A[4][0][50]    = S_in[306];
   assign A[0][1][50]    = S_in[370];
   assign A[1][1][50]    = S_in[434];
   assign A[2][1][50]    = S_in[498];
   assign A[3][1][50]    = S_in[562];
   assign A[4][1][50]    = S_in[626];
   assign A[0][2][50]    = S_in[690];
   assign A[1][2][50]    = S_in[754];
   assign A[2][2][50]    = S_in[818];
   assign A[3][2][50]    = S_in[882];
   assign A[4][2][50]    = S_in[946];
   assign A[0][3][50]    = S_in[1010];
   assign A[1][3][50]    = S_in[1074];
   assign A[2][3][50]    = S_in[1138];
   assign A[3][3][50]    = S_in[1202];
   assign A[4][3][50]    = S_in[1266];
   assign A[0][4][50]    = S_in[1330];
   assign A[1][4][50]    = S_in[1394];
   assign A[2][4][50]    = S_in[1458];
   assign A[3][4][50]    = S_in[1522];
   assign A[4][4][50]    = S_in[1586];
   assign A[0][0][51]    = S_in[51];
   assign A[1][0][51]    = S_in[115];
   assign A[2][0][51]    = S_in[179];
   assign A[3][0][51]    = S_in[243];
   assign A[4][0][51]    = S_in[307];
   assign A[0][1][51]    = S_in[371];
   assign A[1][1][51]    = S_in[435];
   assign A[2][1][51]    = S_in[499];
   assign A[3][1][51]    = S_in[563];
   assign A[4][1][51]    = S_in[627];
   assign A[0][2][51]    = S_in[691];
   assign A[1][2][51]    = S_in[755];
   assign A[2][2][51]    = S_in[819];
   assign A[3][2][51]    = S_in[883];
   assign A[4][2][51]    = S_in[947];
   assign A[0][3][51]    = S_in[1011];
   assign A[1][3][51]    = S_in[1075];
   assign A[2][3][51]    = S_in[1139];
   assign A[3][3][51]    = S_in[1203];
   assign A[4][3][51]    = S_in[1267];
   assign A[0][4][51]    = S_in[1331];
   assign A[1][4][51]    = S_in[1395];
   assign A[2][4][51]    = S_in[1459];
   assign A[3][4][51]    = S_in[1523];
   assign A[4][4][51]    = S_in[1587];
   assign A[0][0][52]    = S_in[52];
   assign A[1][0][52]    = S_in[116];
   assign A[2][0][52]    = S_in[180];
   assign A[3][0][52]    = S_in[244];
   assign A[4][0][52]    = S_in[308];
   assign A[0][1][52]    = S_in[372];
   assign A[1][1][52]    = S_in[436];
   assign A[2][1][52]    = S_in[500];
   assign A[3][1][52]    = S_in[564];
   assign A[4][1][52]    = S_in[628];
   assign A[0][2][52]    = S_in[692];
   assign A[1][2][52]    = S_in[756];
   assign A[2][2][52]    = S_in[820];
   assign A[3][2][52]    = S_in[884];
   assign A[4][2][52]    = S_in[948];
   assign A[0][3][52]    = S_in[1012];
   assign A[1][3][52]    = S_in[1076];
   assign A[2][3][52]    = S_in[1140];
   assign A[3][3][52]    = S_in[1204];
   assign A[4][3][52]    = S_in[1268];
   assign A[0][4][52]    = S_in[1332];
   assign A[1][4][52]    = S_in[1396];
   assign A[2][4][52]    = S_in[1460];
   assign A[3][4][52]    = S_in[1524];
   assign A[4][4][52]    = S_in[1588];
   assign A[0][0][53]    = S_in[53];
   assign A[1][0][53]    = S_in[117];
   assign A[2][0][53]    = S_in[181];
   assign A[3][0][53]    = S_in[245];
   assign A[4][0][53]    = S_in[309];
   assign A[0][1][53]    = S_in[373];
   assign A[1][1][53]    = S_in[437];
   assign A[2][1][53]    = S_in[501];
   assign A[3][1][53]    = S_in[565];
   assign A[4][1][53]    = S_in[629];
   assign A[0][2][53]    = S_in[693];
   assign A[1][2][53]    = S_in[757];
   assign A[2][2][53]    = S_in[821];
   assign A[3][2][53]    = S_in[885];
   assign A[4][2][53]    = S_in[949];
   assign A[0][3][53]    = S_in[1013];
   assign A[1][3][53]    = S_in[1077];
   assign A[2][3][53]    = S_in[1141];
   assign A[3][3][53]    = S_in[1205];
   assign A[4][3][53]    = S_in[1269];
   assign A[0][4][53]    = S_in[1333];
   assign A[1][4][53]    = S_in[1397];
   assign A[2][4][53]    = S_in[1461];
   assign A[3][4][53]    = S_in[1525];
   assign A[4][4][53]    = S_in[1589];
   assign A[0][0][54]    = S_in[54];
   assign A[1][0][54]    = S_in[118];
   assign A[2][0][54]    = S_in[182];
   assign A[3][0][54]    = S_in[246];
   assign A[4][0][54]    = S_in[310];
   assign A[0][1][54]    = S_in[374];
   assign A[1][1][54]    = S_in[438];
   assign A[2][1][54]    = S_in[502];
   assign A[3][1][54]    = S_in[566];
   assign A[4][1][54]    = S_in[630];
   assign A[0][2][54]    = S_in[694];
   assign A[1][2][54]    = S_in[758];
   assign A[2][2][54]    = S_in[822];
   assign A[3][2][54]    = S_in[886];
   assign A[4][2][54]    = S_in[950];
   assign A[0][3][54]    = S_in[1014];
   assign A[1][3][54]    = S_in[1078];
   assign A[2][3][54]    = S_in[1142];
   assign A[3][3][54]    = S_in[1206];
   assign A[4][3][54]    = S_in[1270];
   assign A[0][4][54]    = S_in[1334];
   assign A[1][4][54]    = S_in[1398];
   assign A[2][4][54]    = S_in[1462];
   assign A[3][4][54]    = S_in[1526];
   assign A[4][4][54]    = S_in[1590];
   assign A[0][0][55]    = S_in[55];
   assign A[1][0][55]    = S_in[119];
   assign A[2][0][55]    = S_in[183];
   assign A[3][0][55]    = S_in[247];
   assign A[4][0][55]    = S_in[311];
   assign A[0][1][55]    = S_in[375];
   assign A[1][1][55]    = S_in[439];
   assign A[2][1][55]    = S_in[503];
   assign A[3][1][55]    = S_in[567];
   assign A[4][1][55]    = S_in[631];
   assign A[0][2][55]    = S_in[695];
   assign A[1][2][55]    = S_in[759];
   assign A[2][2][55]    = S_in[823];
   assign A[3][2][55]    = S_in[887];
   assign A[4][2][55]    = S_in[951];
   assign A[0][3][55]    = S_in[1015];
   assign A[1][3][55]    = S_in[1079];
   assign A[2][3][55]    = S_in[1143];
   assign A[3][3][55]    = S_in[1207];
   assign A[4][3][55]    = S_in[1271];
   assign A[0][4][55]    = S_in[1335];
   assign A[1][4][55]    = S_in[1399];
   assign A[2][4][55]    = S_in[1463];
   assign A[3][4][55]    = S_in[1527];
   assign A[4][4][55]    = S_in[1591];
   assign A[0][0][56]    = S_in[56];
   assign A[1][0][56]    = S_in[120];
   assign A[2][0][56]    = S_in[184];
   assign A[3][0][56]    = S_in[248];
   assign A[4][0][56]    = S_in[312];
   assign A[0][1][56]    = S_in[376];
   assign A[1][1][56]    = S_in[440];
   assign A[2][1][56]    = S_in[504];
   assign A[3][1][56]    = S_in[568];
   assign A[4][1][56]    = S_in[632];
   assign A[0][2][56]    = S_in[696];
   assign A[1][2][56]    = S_in[760];
   assign A[2][2][56]    = S_in[824];
   assign A[3][2][56]    = S_in[888];
   assign A[4][2][56]    = S_in[952];
   assign A[0][3][56]    = S_in[1016];
   assign A[1][3][56]    = S_in[1080];
   assign A[2][3][56]    = S_in[1144];
   assign A[3][3][56]    = S_in[1208];
   assign A[4][3][56]    = S_in[1272];
   assign A[0][4][56]    = S_in[1336];
   assign A[1][4][56]    = S_in[1400];
   assign A[2][4][56]    = S_in[1464];
   assign A[3][4][56]    = S_in[1528];
   assign A[4][4][56]    = S_in[1592];
   assign A[0][0][57]    = S_in[57];
   assign A[1][0][57]    = S_in[121];
   assign A[2][0][57]    = S_in[185];
   assign A[3][0][57]    = S_in[249];
   assign A[4][0][57]    = S_in[313];
   assign A[0][1][57]    = S_in[377];
   assign A[1][1][57]    = S_in[441];
   assign A[2][1][57]    = S_in[505];
   assign A[3][1][57]    = S_in[569];
   assign A[4][1][57]    = S_in[633];
   assign A[0][2][57]    = S_in[697];
   assign A[1][2][57]    = S_in[761];
   assign A[2][2][57]    = S_in[825];
   assign A[3][2][57]    = S_in[889];
   assign A[4][2][57]    = S_in[953];
   assign A[0][3][57]    = S_in[1017];
   assign A[1][3][57]    = S_in[1081];
   assign A[2][3][57]    = S_in[1145];
   assign A[3][3][57]    = S_in[1209];
   assign A[4][3][57]    = S_in[1273];
   assign A[0][4][57]    = S_in[1337];
   assign A[1][4][57]    = S_in[1401];
   assign A[2][4][57]    = S_in[1465];
   assign A[3][4][57]    = S_in[1529];
   assign A[4][4][57]    = S_in[1593];
   assign A[0][0][58]    = S_in[58];
   assign A[1][0][58]    = S_in[122];
   assign A[2][0][58]    = S_in[186];
   assign A[3][0][58]    = S_in[250];
   assign A[4][0][58]    = S_in[314];
   assign A[0][1][58]    = S_in[378];
   assign A[1][1][58]    = S_in[442];
   assign A[2][1][58]    = S_in[506];
   assign A[3][1][58]    = S_in[570];
   assign A[4][1][58]    = S_in[634];
   assign A[0][2][58]    = S_in[698];
   assign A[1][2][58]    = S_in[762];
   assign A[2][2][58]    = S_in[826];
   assign A[3][2][58]    = S_in[890];
   assign A[4][2][58]    = S_in[954];
   assign A[0][3][58]    = S_in[1018];
   assign A[1][3][58]    = S_in[1082];
   assign A[2][3][58]    = S_in[1146];
   assign A[3][3][58]    = S_in[1210];
   assign A[4][3][58]    = S_in[1274];
   assign A[0][4][58]    = S_in[1338];
   assign A[1][4][58]    = S_in[1402];
   assign A[2][4][58]    = S_in[1466];
   assign A[3][4][58]    = S_in[1530];
   assign A[4][4][58]    = S_in[1594];
   assign A[0][0][59]    = S_in[59];
   assign A[1][0][59]    = S_in[123];
   assign A[2][0][59]    = S_in[187];
   assign A[3][0][59]    = S_in[251];
   assign A[4][0][59]    = S_in[315];
   assign A[0][1][59]    = S_in[379];
   assign A[1][1][59]    = S_in[443];
   assign A[2][1][59]    = S_in[507];
   assign A[3][1][59]    = S_in[571];
   assign A[4][1][59]    = S_in[635];
   assign A[0][2][59]    = S_in[699];
   assign A[1][2][59]    = S_in[763];
   assign A[2][2][59]    = S_in[827];
   assign A[3][2][59]    = S_in[891];
   assign A[4][2][59]    = S_in[955];
   assign A[0][3][59]    = S_in[1019];
   assign A[1][3][59]    = S_in[1083];
   assign A[2][3][59]    = S_in[1147];
   assign A[3][3][59]    = S_in[1211];
   assign A[4][3][59]    = S_in[1275];
   assign A[0][4][59]    = S_in[1339];
   assign A[1][4][59]    = S_in[1403];
   assign A[2][4][59]    = S_in[1467];
   assign A[3][4][59]    = S_in[1531];
   assign A[4][4][59]    = S_in[1595];
   assign A[0][0][60]    = S_in[60];
   assign A[1][0][60]    = S_in[124];
   assign A[2][0][60]    = S_in[188];
   assign A[3][0][60]    = S_in[252];
   assign A[4][0][60]    = S_in[316];
   assign A[0][1][60]    = S_in[380];
   assign A[1][1][60]    = S_in[444];
   assign A[2][1][60]    = S_in[508];
   assign A[3][1][60]    = S_in[572];
   assign A[4][1][60]    = S_in[636];
   assign A[0][2][60]    = S_in[700];
   assign A[1][2][60]    = S_in[764];
   assign A[2][2][60]    = S_in[828];
   assign A[3][2][60]    = S_in[892];
   assign A[4][2][60]    = S_in[956];
   assign A[0][3][60]    = S_in[1020];
   assign A[1][3][60]    = S_in[1084];
   assign A[2][3][60]    = S_in[1148];
   assign A[3][3][60]    = S_in[1212];
   assign A[4][3][60]    = S_in[1276];
   assign A[0][4][60]    = S_in[1340];
   assign A[1][4][60]    = S_in[1404];
   assign A[2][4][60]    = S_in[1468];
   assign A[3][4][60]    = S_in[1532];
   assign A[4][4][60]    = S_in[1596];
   assign A[0][0][61]    = S_in[61];
   assign A[1][0][61]    = S_in[125];
   assign A[2][0][61]    = S_in[189];
   assign A[3][0][61]    = S_in[253];
   assign A[4][0][61]    = S_in[317];
   assign A[0][1][61]    = S_in[381];
   assign A[1][1][61]    = S_in[445];
   assign A[2][1][61]    = S_in[509];
   assign A[3][1][61]    = S_in[573];
   assign A[4][1][61]    = S_in[637];
   assign A[0][2][61]    = S_in[701];
   assign A[1][2][61]    = S_in[765];
   assign A[2][2][61]    = S_in[829];
   assign A[3][2][61]    = S_in[893];
   assign A[4][2][61]    = S_in[957];
   assign A[0][3][61]    = S_in[1021];
   assign A[1][3][61]    = S_in[1085];
   assign A[2][3][61]    = S_in[1149];
   assign A[3][3][61]    = S_in[1213];
   assign A[4][3][61]    = S_in[1277];
   assign A[0][4][61]    = S_in[1341];
   assign A[1][4][61]    = S_in[1405];
   assign A[2][4][61]    = S_in[1469];
   assign A[3][4][61]    = S_in[1533];
   assign A[4][4][61]    = S_in[1597];
   assign A[0][0][62]    = S_in[62];
   assign A[1][0][62]    = S_in[126];
   assign A[2][0][62]    = S_in[190];
   assign A[3][0][62]    = S_in[254];
   assign A[4][0][62]    = S_in[318];
   assign A[0][1][62]    = S_in[382];
   assign A[1][1][62]    = S_in[446];
   assign A[2][1][62]    = S_in[510];
   assign A[3][1][62]    = S_in[574];
   assign A[4][1][62]    = S_in[638];
   assign A[0][2][62]    = S_in[702];
   assign A[1][2][62]    = S_in[766];
   assign A[2][2][62]    = S_in[830];
   assign A[3][2][62]    = S_in[894];
   assign A[4][2][62]    = S_in[958];
   assign A[0][3][62]    = S_in[1022];
   assign A[1][3][62]    = S_in[1086];
   assign A[2][3][62]    = S_in[1150];
   assign A[3][3][62]    = S_in[1214];
   assign A[4][3][62]    = S_in[1278];
   assign A[0][4][62]    = S_in[1342];
   assign A[1][4][62]    = S_in[1406];
   assign A[2][4][62]    = S_in[1470];
   assign A[3][4][62]    = S_in[1534];
   assign A[4][4][62]    = S_in[1598];
   assign A[0][0][63]    = S_in[63];
   assign A[1][0][63]    = S_in[127];
   assign A[2][0][63]    = S_in[191];
   assign A[3][0][63]    = S_in[255];
   assign A[4][0][63]    = S_in[319];
   assign A[0][1][63]    = S_in[383];
   assign A[1][1][63]    = S_in[447];
   assign A[2][1][63]    = S_in[511];
   assign A[3][1][63]    = S_in[575];
   assign A[4][1][63]    = S_in[639];
   assign A[0][2][63]    = S_in[703];
   assign A[1][2][63]    = S_in[767];
   assign A[2][2][63]    = S_in[831];
   assign A[3][2][63]    = S_in[895];
   assign A[4][2][63]    = S_in[959];
   assign A[0][3][63]    = S_in[1023];
   assign A[1][3][63]    = S_in[1087];
   assign A[2][3][63]    = S_in[1151];
   assign A[3][3][63]    = S_in[1215];
   assign A[4][3][63]    = S_in[1279];
   assign A[0][4][63]    = S_in[1343];
   assign A[1][4][63]    = S_in[1407];
   assign A[2][4][63]    = S_in[1471];
   assign A[3][4][63]    = S_in[1535];
   assign A[4][4][63]    = S_in[1599];
//--------------------------- THETA ---------------------------
    // Step 1: Compute C[x][z]
    assign C[0][0]     = A[0][0][0] ^ A[0][1][0] ^ A[0][2][0] ^ A[0][3][0] ^ A[0][4][0];
    assign C[0][1]     = A[0][0][1] ^ A[0][1][1] ^ A[0][2][1] ^ A[0][3][1] ^ A[0][4][1];
    assign C[0][2]     = A[0][0][2] ^ A[0][1][2] ^ A[0][2][2] ^ A[0][3][2] ^ A[0][4][2];
    assign C[0][3]     = A[0][0][3] ^ A[0][1][3] ^ A[0][2][3] ^ A[0][3][3] ^ A[0][4][3];
    assign C[0][4]     = A[0][0][4] ^ A[0][1][4] ^ A[0][2][4] ^ A[0][3][4] ^ A[0][4][4];
    assign C[0][5]     = A[0][0][5] ^ A[0][1][5] ^ A[0][2][5] ^ A[0][3][5] ^ A[0][4][5];
    assign C[0][6]     = A[0][0][6] ^ A[0][1][6] ^ A[0][2][6] ^ A[0][3][6] ^ A[0][4][6];
    assign C[0][7]     = A[0][0][7] ^ A[0][1][7] ^ A[0][2][7] ^ A[0][3][7] ^ A[0][4][7];
    assign C[0][8]     = A[0][0][8] ^ A[0][1][8] ^ A[0][2][8] ^ A[0][3][8] ^ A[0][4][8];
    assign C[0][9]     = A[0][0][9] ^ A[0][1][9] ^ A[0][2][9] ^ A[0][3][9] ^ A[0][4][9];
    assign C[0][10]     = A[0][0][10] ^ A[0][1][10] ^ A[0][2][10] ^ A[0][3][10] ^ A[0][4][10];
    assign C[0][11]     = A[0][0][11] ^ A[0][1][11] ^ A[0][2][11] ^ A[0][3][11] ^ A[0][4][11];
    assign C[0][12]     = A[0][0][12] ^ A[0][1][12] ^ A[0][2][12] ^ A[0][3][12] ^ A[0][4][12];
    assign C[0][13]     = A[0][0][13] ^ A[0][1][13] ^ A[0][2][13] ^ A[0][3][13] ^ A[0][4][13];
    assign C[0][14]     = A[0][0][14] ^ A[0][1][14] ^ A[0][2][14] ^ A[0][3][14] ^ A[0][4][14];
    assign C[0][15]     = A[0][0][15] ^ A[0][1][15] ^ A[0][2][15] ^ A[0][3][15] ^ A[0][4][15];
    assign C[0][16]     = A[0][0][16] ^ A[0][1][16] ^ A[0][2][16] ^ A[0][3][16] ^ A[0][4][16];
    assign C[0][17]     = A[0][0][17] ^ A[0][1][17] ^ A[0][2][17] ^ A[0][3][17] ^ A[0][4][17];
    assign C[0][18]     = A[0][0][18] ^ A[0][1][18] ^ A[0][2][18] ^ A[0][3][18] ^ A[0][4][18];
    assign C[0][19]     = A[0][0][19] ^ A[0][1][19] ^ A[0][2][19] ^ A[0][3][19] ^ A[0][4][19];
    assign C[0][20]     = A[0][0][20] ^ A[0][1][20] ^ A[0][2][20] ^ A[0][3][20] ^ A[0][4][20];
    assign C[0][21]     = A[0][0][21] ^ A[0][1][21] ^ A[0][2][21] ^ A[0][3][21] ^ A[0][4][21];
    assign C[0][22]     = A[0][0][22] ^ A[0][1][22] ^ A[0][2][22] ^ A[0][3][22] ^ A[0][4][22];
    assign C[0][23]     = A[0][0][23] ^ A[0][1][23] ^ A[0][2][23] ^ A[0][3][23] ^ A[0][4][23];
    assign C[0][24]     = A[0][0][24] ^ A[0][1][24] ^ A[0][2][24] ^ A[0][3][24] ^ A[0][4][24];
    assign C[0][25]     = A[0][0][25] ^ A[0][1][25] ^ A[0][2][25] ^ A[0][3][25] ^ A[0][4][25];
    assign C[0][26]     = A[0][0][26] ^ A[0][1][26] ^ A[0][2][26] ^ A[0][3][26] ^ A[0][4][26];
    assign C[0][27]     = A[0][0][27] ^ A[0][1][27] ^ A[0][2][27] ^ A[0][3][27] ^ A[0][4][27];
    assign C[0][28]     = A[0][0][28] ^ A[0][1][28] ^ A[0][2][28] ^ A[0][3][28] ^ A[0][4][28];
    assign C[0][29]     = A[0][0][29] ^ A[0][1][29] ^ A[0][2][29] ^ A[0][3][29] ^ A[0][4][29];
    assign C[0][30]     = A[0][0][30] ^ A[0][1][30] ^ A[0][2][30] ^ A[0][3][30] ^ A[0][4][30];
    assign C[0][31]     = A[0][0][31] ^ A[0][1][31] ^ A[0][2][31] ^ A[0][3][31] ^ A[0][4][31];
    assign C[0][32]     = A[0][0][32] ^ A[0][1][32] ^ A[0][2][32] ^ A[0][3][32] ^ A[0][4][32];
    assign C[0][33]     = A[0][0][33] ^ A[0][1][33] ^ A[0][2][33] ^ A[0][3][33] ^ A[0][4][33];
    assign C[0][34]     = A[0][0][34] ^ A[0][1][34] ^ A[0][2][34] ^ A[0][3][34] ^ A[0][4][34];
    assign C[0][35]     = A[0][0][35] ^ A[0][1][35] ^ A[0][2][35] ^ A[0][3][35] ^ A[0][4][35];
    assign C[0][36]     = A[0][0][36] ^ A[0][1][36] ^ A[0][2][36] ^ A[0][3][36] ^ A[0][4][36];
    assign C[0][37]     = A[0][0][37] ^ A[0][1][37] ^ A[0][2][37] ^ A[0][3][37] ^ A[0][4][37];
    assign C[0][38]     = A[0][0][38] ^ A[0][1][38] ^ A[0][2][38] ^ A[0][3][38] ^ A[0][4][38];
    assign C[0][39]     = A[0][0][39] ^ A[0][1][39] ^ A[0][2][39] ^ A[0][3][39] ^ A[0][4][39];
    assign C[0][40]     = A[0][0][40] ^ A[0][1][40] ^ A[0][2][40] ^ A[0][3][40] ^ A[0][4][40];
    assign C[0][41]     = A[0][0][41] ^ A[0][1][41] ^ A[0][2][41] ^ A[0][3][41] ^ A[0][4][41];
    assign C[0][42]     = A[0][0][42] ^ A[0][1][42] ^ A[0][2][42] ^ A[0][3][42] ^ A[0][4][42];
    assign C[0][43]     = A[0][0][43] ^ A[0][1][43] ^ A[0][2][43] ^ A[0][3][43] ^ A[0][4][43];
    assign C[0][44]     = A[0][0][44] ^ A[0][1][44] ^ A[0][2][44] ^ A[0][3][44] ^ A[0][4][44];
    assign C[0][45]     = A[0][0][45] ^ A[0][1][45] ^ A[0][2][45] ^ A[0][3][45] ^ A[0][4][45];
    assign C[0][46]     = A[0][0][46] ^ A[0][1][46] ^ A[0][2][46] ^ A[0][3][46] ^ A[0][4][46];
    assign C[0][47]     = A[0][0][47] ^ A[0][1][47] ^ A[0][2][47] ^ A[0][3][47] ^ A[0][4][47];
    assign C[0][48]     = A[0][0][48] ^ A[0][1][48] ^ A[0][2][48] ^ A[0][3][48] ^ A[0][4][48];
    assign C[0][49]     = A[0][0][49] ^ A[0][1][49] ^ A[0][2][49] ^ A[0][3][49] ^ A[0][4][49];
    assign C[0][50]     = A[0][0][50] ^ A[0][1][50] ^ A[0][2][50] ^ A[0][3][50] ^ A[0][4][50];
    assign C[0][51]     = A[0][0][51] ^ A[0][1][51] ^ A[0][2][51] ^ A[0][3][51] ^ A[0][4][51];
    assign C[0][52]     = A[0][0][52] ^ A[0][1][52] ^ A[0][2][52] ^ A[0][3][52] ^ A[0][4][52];
    assign C[0][53]     = A[0][0][53] ^ A[0][1][53] ^ A[0][2][53] ^ A[0][3][53] ^ A[0][4][53];
    assign C[0][54]     = A[0][0][54] ^ A[0][1][54] ^ A[0][2][54] ^ A[0][3][54] ^ A[0][4][54];
    assign C[0][55]     = A[0][0][55] ^ A[0][1][55] ^ A[0][2][55] ^ A[0][3][55] ^ A[0][4][55];
    assign C[0][56]     = A[0][0][56] ^ A[0][1][56] ^ A[0][2][56] ^ A[0][3][56] ^ A[0][4][56];
    assign C[0][57]     = A[0][0][57] ^ A[0][1][57] ^ A[0][2][57] ^ A[0][3][57] ^ A[0][4][57];
    assign C[0][58]     = A[0][0][58] ^ A[0][1][58] ^ A[0][2][58] ^ A[0][3][58] ^ A[0][4][58];
    assign C[0][59]     = A[0][0][59] ^ A[0][1][59] ^ A[0][2][59] ^ A[0][3][59] ^ A[0][4][59];
    assign C[0][60]     = A[0][0][60] ^ A[0][1][60] ^ A[0][2][60] ^ A[0][3][60] ^ A[0][4][60];
    assign C[0][61]     = A[0][0][61] ^ A[0][1][61] ^ A[0][2][61] ^ A[0][3][61] ^ A[0][4][61];
    assign C[0][62]     = A[0][0][62] ^ A[0][1][62] ^ A[0][2][62] ^ A[0][3][62] ^ A[0][4][62];
    assign C[0][63]     = A[0][0][63] ^ A[0][1][63] ^ A[0][2][63] ^ A[0][3][63] ^ A[0][4][63];
    assign C[1][0]     = A[1][0][0] ^ A[1][1][0] ^ A[1][2][0] ^ A[1][3][0] ^ A[1][4][0];
    assign C[1][1]     = A[1][0][1] ^ A[1][1][1] ^ A[1][2][1] ^ A[1][3][1] ^ A[1][4][1];
    assign C[1][2]     = A[1][0][2] ^ A[1][1][2] ^ A[1][2][2] ^ A[1][3][2] ^ A[1][4][2];
    assign C[1][3]     = A[1][0][3] ^ A[1][1][3] ^ A[1][2][3] ^ A[1][3][3] ^ A[1][4][3];
    assign C[1][4]     = A[1][0][4] ^ A[1][1][4] ^ A[1][2][4] ^ A[1][3][4] ^ A[1][4][4];
    assign C[1][5]     = A[1][0][5] ^ A[1][1][5] ^ A[1][2][5] ^ A[1][3][5] ^ A[1][4][5];
    assign C[1][6]     = A[1][0][6] ^ A[1][1][6] ^ A[1][2][6] ^ A[1][3][6] ^ A[1][4][6];
    assign C[1][7]     = A[1][0][7] ^ A[1][1][7] ^ A[1][2][7] ^ A[1][3][7] ^ A[1][4][7];
    assign C[1][8]     = A[1][0][8] ^ A[1][1][8] ^ A[1][2][8] ^ A[1][3][8] ^ A[1][4][8];
    assign C[1][9]     = A[1][0][9] ^ A[1][1][9] ^ A[1][2][9] ^ A[1][3][9] ^ A[1][4][9];
    assign C[1][10]     = A[1][0][10] ^ A[1][1][10] ^ A[1][2][10] ^ A[1][3][10] ^ A[1][4][10];
    assign C[1][11]     = A[1][0][11] ^ A[1][1][11] ^ A[1][2][11] ^ A[1][3][11] ^ A[1][4][11];
    assign C[1][12]     = A[1][0][12] ^ A[1][1][12] ^ A[1][2][12] ^ A[1][3][12] ^ A[1][4][12];
    assign C[1][13]     = A[1][0][13] ^ A[1][1][13] ^ A[1][2][13] ^ A[1][3][13] ^ A[1][4][13];
    assign C[1][14]     = A[1][0][14] ^ A[1][1][14] ^ A[1][2][14] ^ A[1][3][14] ^ A[1][4][14];
    assign C[1][15]     = A[1][0][15] ^ A[1][1][15] ^ A[1][2][15] ^ A[1][3][15] ^ A[1][4][15];
    assign C[1][16]     = A[1][0][16] ^ A[1][1][16] ^ A[1][2][16] ^ A[1][3][16] ^ A[1][4][16];
    assign C[1][17]     = A[1][0][17] ^ A[1][1][17] ^ A[1][2][17] ^ A[1][3][17] ^ A[1][4][17];
    assign C[1][18]     = A[1][0][18] ^ A[1][1][18] ^ A[1][2][18] ^ A[1][3][18] ^ A[1][4][18];
    assign C[1][19]     = A[1][0][19] ^ A[1][1][19] ^ A[1][2][19] ^ A[1][3][19] ^ A[1][4][19];
    assign C[1][20]     = A[1][0][20] ^ A[1][1][20] ^ A[1][2][20] ^ A[1][3][20] ^ A[1][4][20];
    assign C[1][21]     = A[1][0][21] ^ A[1][1][21] ^ A[1][2][21] ^ A[1][3][21] ^ A[1][4][21];
    assign C[1][22]     = A[1][0][22] ^ A[1][1][22] ^ A[1][2][22] ^ A[1][3][22] ^ A[1][4][22];
    assign C[1][23]     = A[1][0][23] ^ A[1][1][23] ^ A[1][2][23] ^ A[1][3][23] ^ A[1][4][23];
    assign C[1][24]     = A[1][0][24] ^ A[1][1][24] ^ A[1][2][24] ^ A[1][3][24] ^ A[1][4][24];
    assign C[1][25]     = A[1][0][25] ^ A[1][1][25] ^ A[1][2][25] ^ A[1][3][25] ^ A[1][4][25];
    assign C[1][26]     = A[1][0][26] ^ A[1][1][26] ^ A[1][2][26] ^ A[1][3][26] ^ A[1][4][26];
    assign C[1][27]     = A[1][0][27] ^ A[1][1][27] ^ A[1][2][27] ^ A[1][3][27] ^ A[1][4][27];
    assign C[1][28]     = A[1][0][28] ^ A[1][1][28] ^ A[1][2][28] ^ A[1][3][28] ^ A[1][4][28];
    assign C[1][29]     = A[1][0][29] ^ A[1][1][29] ^ A[1][2][29] ^ A[1][3][29] ^ A[1][4][29];
    assign C[1][30]     = A[1][0][30] ^ A[1][1][30] ^ A[1][2][30] ^ A[1][3][30] ^ A[1][4][30];
    assign C[1][31]     = A[1][0][31] ^ A[1][1][31] ^ A[1][2][31] ^ A[1][3][31] ^ A[1][4][31];
    assign C[1][32]     = A[1][0][32] ^ A[1][1][32] ^ A[1][2][32] ^ A[1][3][32] ^ A[1][4][32];
    assign C[1][33]     = A[1][0][33] ^ A[1][1][33] ^ A[1][2][33] ^ A[1][3][33] ^ A[1][4][33];
    assign C[1][34]     = A[1][0][34] ^ A[1][1][34] ^ A[1][2][34] ^ A[1][3][34] ^ A[1][4][34];
    assign C[1][35]     = A[1][0][35] ^ A[1][1][35] ^ A[1][2][35] ^ A[1][3][35] ^ A[1][4][35];
    assign C[1][36]     = A[1][0][36] ^ A[1][1][36] ^ A[1][2][36] ^ A[1][3][36] ^ A[1][4][36];
    assign C[1][37]     = A[1][0][37] ^ A[1][1][37] ^ A[1][2][37] ^ A[1][3][37] ^ A[1][4][37];
    assign C[1][38]     = A[1][0][38] ^ A[1][1][38] ^ A[1][2][38] ^ A[1][3][38] ^ A[1][4][38];
    assign C[1][39]     = A[1][0][39] ^ A[1][1][39] ^ A[1][2][39] ^ A[1][3][39] ^ A[1][4][39];
    assign C[1][40]     = A[1][0][40] ^ A[1][1][40] ^ A[1][2][40] ^ A[1][3][40] ^ A[1][4][40];
    assign C[1][41]     = A[1][0][41] ^ A[1][1][41] ^ A[1][2][41] ^ A[1][3][41] ^ A[1][4][41];
    assign C[1][42]     = A[1][0][42] ^ A[1][1][42] ^ A[1][2][42] ^ A[1][3][42] ^ A[1][4][42];
    assign C[1][43]     = A[1][0][43] ^ A[1][1][43] ^ A[1][2][43] ^ A[1][3][43] ^ A[1][4][43];
    assign C[1][44]     = A[1][0][44] ^ A[1][1][44] ^ A[1][2][44] ^ A[1][3][44] ^ A[1][4][44];
    assign C[1][45]     = A[1][0][45] ^ A[1][1][45] ^ A[1][2][45] ^ A[1][3][45] ^ A[1][4][45];
    assign C[1][46]     = A[1][0][46] ^ A[1][1][46] ^ A[1][2][46] ^ A[1][3][46] ^ A[1][4][46];
    assign C[1][47]     = A[1][0][47] ^ A[1][1][47] ^ A[1][2][47] ^ A[1][3][47] ^ A[1][4][47];
    assign C[1][48]     = A[1][0][48] ^ A[1][1][48] ^ A[1][2][48] ^ A[1][3][48] ^ A[1][4][48];
    assign C[1][49]     = A[1][0][49] ^ A[1][1][49] ^ A[1][2][49] ^ A[1][3][49] ^ A[1][4][49];
    assign C[1][50]     = A[1][0][50] ^ A[1][1][50] ^ A[1][2][50] ^ A[1][3][50] ^ A[1][4][50];
    assign C[1][51]     = A[1][0][51] ^ A[1][1][51] ^ A[1][2][51] ^ A[1][3][51] ^ A[1][4][51];
    assign C[1][52]     = A[1][0][52] ^ A[1][1][52] ^ A[1][2][52] ^ A[1][3][52] ^ A[1][4][52];
    assign C[1][53]     = A[1][0][53] ^ A[1][1][53] ^ A[1][2][53] ^ A[1][3][53] ^ A[1][4][53];
    assign C[1][54]     = A[1][0][54] ^ A[1][1][54] ^ A[1][2][54] ^ A[1][3][54] ^ A[1][4][54];
    assign C[1][55]     = A[1][0][55] ^ A[1][1][55] ^ A[1][2][55] ^ A[1][3][55] ^ A[1][4][55];
    assign C[1][56]     = A[1][0][56] ^ A[1][1][56] ^ A[1][2][56] ^ A[1][3][56] ^ A[1][4][56];
    assign C[1][57]     = A[1][0][57] ^ A[1][1][57] ^ A[1][2][57] ^ A[1][3][57] ^ A[1][4][57];
    assign C[1][58]     = A[1][0][58] ^ A[1][1][58] ^ A[1][2][58] ^ A[1][3][58] ^ A[1][4][58];
    assign C[1][59]     = A[1][0][59] ^ A[1][1][59] ^ A[1][2][59] ^ A[1][3][59] ^ A[1][4][59];
    assign C[1][60]     = A[1][0][60] ^ A[1][1][60] ^ A[1][2][60] ^ A[1][3][60] ^ A[1][4][60];
    assign C[1][61]     = A[1][0][61] ^ A[1][1][61] ^ A[1][2][61] ^ A[1][3][61] ^ A[1][4][61];
    assign C[1][62]     = A[1][0][62] ^ A[1][1][62] ^ A[1][2][62] ^ A[1][3][62] ^ A[1][4][62];
    assign C[1][63]     = A[1][0][63] ^ A[1][1][63] ^ A[1][2][63] ^ A[1][3][63] ^ A[1][4][63];
    assign C[2][0]     = A[2][0][0] ^ A[2][1][0] ^ A[2][2][0] ^ A[2][3][0] ^ A[2][4][0];
    assign C[2][1]     = A[2][0][1] ^ A[2][1][1] ^ A[2][2][1] ^ A[2][3][1] ^ A[2][4][1];
    assign C[2][2]     = A[2][0][2] ^ A[2][1][2] ^ A[2][2][2] ^ A[2][3][2] ^ A[2][4][2];
    assign C[2][3]     = A[2][0][3] ^ A[2][1][3] ^ A[2][2][3] ^ A[2][3][3] ^ A[2][4][3];
    assign C[2][4]     = A[2][0][4] ^ A[2][1][4] ^ A[2][2][4] ^ A[2][3][4] ^ A[2][4][4];
    assign C[2][5]     = A[2][0][5] ^ A[2][1][5] ^ A[2][2][5] ^ A[2][3][5] ^ A[2][4][5];
    assign C[2][6]     = A[2][0][6] ^ A[2][1][6] ^ A[2][2][6] ^ A[2][3][6] ^ A[2][4][6];
    assign C[2][7]     = A[2][0][7] ^ A[2][1][7] ^ A[2][2][7] ^ A[2][3][7] ^ A[2][4][7];
    assign C[2][8]     = A[2][0][8] ^ A[2][1][8] ^ A[2][2][8] ^ A[2][3][8] ^ A[2][4][8];
    assign C[2][9]     = A[2][0][9] ^ A[2][1][9] ^ A[2][2][9] ^ A[2][3][9] ^ A[2][4][9];
    assign C[2][10]     = A[2][0][10] ^ A[2][1][10] ^ A[2][2][10] ^ A[2][3][10] ^ A[2][4][10];
    assign C[2][11]     = A[2][0][11] ^ A[2][1][11] ^ A[2][2][11] ^ A[2][3][11] ^ A[2][4][11];
    assign C[2][12]     = A[2][0][12] ^ A[2][1][12] ^ A[2][2][12] ^ A[2][3][12] ^ A[2][4][12];
    assign C[2][13]     = A[2][0][13] ^ A[2][1][13] ^ A[2][2][13] ^ A[2][3][13] ^ A[2][4][13];
    assign C[2][14]     = A[2][0][14] ^ A[2][1][14] ^ A[2][2][14] ^ A[2][3][14] ^ A[2][4][14];
    assign C[2][15]     = A[2][0][15] ^ A[2][1][15] ^ A[2][2][15] ^ A[2][3][15] ^ A[2][4][15];
    assign C[2][16]     = A[2][0][16] ^ A[2][1][16] ^ A[2][2][16] ^ A[2][3][16] ^ A[2][4][16];
    assign C[2][17]     = A[2][0][17] ^ A[2][1][17] ^ A[2][2][17] ^ A[2][3][17] ^ A[2][4][17];
    assign C[2][18]     = A[2][0][18] ^ A[2][1][18] ^ A[2][2][18] ^ A[2][3][18] ^ A[2][4][18];
    assign C[2][19]     = A[2][0][19] ^ A[2][1][19] ^ A[2][2][19] ^ A[2][3][19] ^ A[2][4][19];
    assign C[2][20]     = A[2][0][20] ^ A[2][1][20] ^ A[2][2][20] ^ A[2][3][20] ^ A[2][4][20];
    assign C[2][21]     = A[2][0][21] ^ A[2][1][21] ^ A[2][2][21] ^ A[2][3][21] ^ A[2][4][21];
    assign C[2][22]     = A[2][0][22] ^ A[2][1][22] ^ A[2][2][22] ^ A[2][3][22] ^ A[2][4][22];
    assign C[2][23]     = A[2][0][23] ^ A[2][1][23] ^ A[2][2][23] ^ A[2][3][23] ^ A[2][4][23];
    assign C[2][24]     = A[2][0][24] ^ A[2][1][24] ^ A[2][2][24] ^ A[2][3][24] ^ A[2][4][24];
    assign C[2][25]     = A[2][0][25] ^ A[2][1][25] ^ A[2][2][25] ^ A[2][3][25] ^ A[2][4][25];
    assign C[2][26]     = A[2][0][26] ^ A[2][1][26] ^ A[2][2][26] ^ A[2][3][26] ^ A[2][4][26];
    assign C[2][27]     = A[2][0][27] ^ A[2][1][27] ^ A[2][2][27] ^ A[2][3][27] ^ A[2][4][27];
    assign C[2][28]     = A[2][0][28] ^ A[2][1][28] ^ A[2][2][28] ^ A[2][3][28] ^ A[2][4][28];
    assign C[2][29]     = A[2][0][29] ^ A[2][1][29] ^ A[2][2][29] ^ A[2][3][29] ^ A[2][4][29];
    assign C[2][30]     = A[2][0][30] ^ A[2][1][30] ^ A[2][2][30] ^ A[2][3][30] ^ A[2][4][30];
    assign C[2][31]     = A[2][0][31] ^ A[2][1][31] ^ A[2][2][31] ^ A[2][3][31] ^ A[2][4][31];
    assign C[2][32]     = A[2][0][32] ^ A[2][1][32] ^ A[2][2][32] ^ A[2][3][32] ^ A[2][4][32];
    assign C[2][33]     = A[2][0][33] ^ A[2][1][33] ^ A[2][2][33] ^ A[2][3][33] ^ A[2][4][33];
    assign C[2][34]     = A[2][0][34] ^ A[2][1][34] ^ A[2][2][34] ^ A[2][3][34] ^ A[2][4][34];
    assign C[2][35]     = A[2][0][35] ^ A[2][1][35] ^ A[2][2][35] ^ A[2][3][35] ^ A[2][4][35];
    assign C[2][36]     = A[2][0][36] ^ A[2][1][36] ^ A[2][2][36] ^ A[2][3][36] ^ A[2][4][36];
    assign C[2][37]     = A[2][0][37] ^ A[2][1][37] ^ A[2][2][37] ^ A[2][3][37] ^ A[2][4][37];
    assign C[2][38]     = A[2][0][38] ^ A[2][1][38] ^ A[2][2][38] ^ A[2][3][38] ^ A[2][4][38];
    assign C[2][39]     = A[2][0][39] ^ A[2][1][39] ^ A[2][2][39] ^ A[2][3][39] ^ A[2][4][39];
    assign C[2][40]     = A[2][0][40] ^ A[2][1][40] ^ A[2][2][40] ^ A[2][3][40] ^ A[2][4][40];
    assign C[2][41]     = A[2][0][41] ^ A[2][1][41] ^ A[2][2][41] ^ A[2][3][41] ^ A[2][4][41];
    assign C[2][42]     = A[2][0][42] ^ A[2][1][42] ^ A[2][2][42] ^ A[2][3][42] ^ A[2][4][42];
    assign C[2][43]     = A[2][0][43] ^ A[2][1][43] ^ A[2][2][43] ^ A[2][3][43] ^ A[2][4][43];
    assign C[2][44]     = A[2][0][44] ^ A[2][1][44] ^ A[2][2][44] ^ A[2][3][44] ^ A[2][4][44];
    assign C[2][45]     = A[2][0][45] ^ A[2][1][45] ^ A[2][2][45] ^ A[2][3][45] ^ A[2][4][45];
    assign C[2][46]     = A[2][0][46] ^ A[2][1][46] ^ A[2][2][46] ^ A[2][3][46] ^ A[2][4][46];
    assign C[2][47]     = A[2][0][47] ^ A[2][1][47] ^ A[2][2][47] ^ A[2][3][47] ^ A[2][4][47];
    assign C[2][48]     = A[2][0][48] ^ A[2][1][48] ^ A[2][2][48] ^ A[2][3][48] ^ A[2][4][48];
    assign C[2][49]     = A[2][0][49] ^ A[2][1][49] ^ A[2][2][49] ^ A[2][3][49] ^ A[2][4][49];
    assign C[2][50]     = A[2][0][50] ^ A[2][1][50] ^ A[2][2][50] ^ A[2][3][50] ^ A[2][4][50];
    assign C[2][51]     = A[2][0][51] ^ A[2][1][51] ^ A[2][2][51] ^ A[2][3][51] ^ A[2][4][51];
    assign C[2][52]     = A[2][0][52] ^ A[2][1][52] ^ A[2][2][52] ^ A[2][3][52] ^ A[2][4][52];
    assign C[2][53]     = A[2][0][53] ^ A[2][1][53] ^ A[2][2][53] ^ A[2][3][53] ^ A[2][4][53];
    assign C[2][54]     = A[2][0][54] ^ A[2][1][54] ^ A[2][2][54] ^ A[2][3][54] ^ A[2][4][54];
    assign C[2][55]     = A[2][0][55] ^ A[2][1][55] ^ A[2][2][55] ^ A[2][3][55] ^ A[2][4][55];
    assign C[2][56]     = A[2][0][56] ^ A[2][1][56] ^ A[2][2][56] ^ A[2][3][56] ^ A[2][4][56];
    assign C[2][57]     = A[2][0][57] ^ A[2][1][57] ^ A[2][2][57] ^ A[2][3][57] ^ A[2][4][57];
    assign C[2][58]     = A[2][0][58] ^ A[2][1][58] ^ A[2][2][58] ^ A[2][3][58] ^ A[2][4][58];
    assign C[2][59]     = A[2][0][59] ^ A[2][1][59] ^ A[2][2][59] ^ A[2][3][59] ^ A[2][4][59];
    assign C[2][60]     = A[2][0][60] ^ A[2][1][60] ^ A[2][2][60] ^ A[2][3][60] ^ A[2][4][60];
    assign C[2][61]     = A[2][0][61] ^ A[2][1][61] ^ A[2][2][61] ^ A[2][3][61] ^ A[2][4][61];
    assign C[2][62]     = A[2][0][62] ^ A[2][1][62] ^ A[2][2][62] ^ A[2][3][62] ^ A[2][4][62];
    assign C[2][63]     = A[2][0][63] ^ A[2][1][63] ^ A[2][2][63] ^ A[2][3][63] ^ A[2][4][63];
    assign C[3][0]     = A[3][0][0] ^ A[3][1][0] ^ A[3][2][0] ^ A[3][3][0] ^ A[3][4][0];
    assign C[3][1]     = A[3][0][1] ^ A[3][1][1] ^ A[3][2][1] ^ A[3][3][1] ^ A[3][4][1];
    assign C[3][2]     = A[3][0][2] ^ A[3][1][2] ^ A[3][2][2] ^ A[3][3][2] ^ A[3][4][2];
    assign C[3][3]     = A[3][0][3] ^ A[3][1][3] ^ A[3][2][3] ^ A[3][3][3] ^ A[3][4][3];
    assign C[3][4]     = A[3][0][4] ^ A[3][1][4] ^ A[3][2][4] ^ A[3][3][4] ^ A[3][4][4];
    assign C[3][5]     = A[3][0][5] ^ A[3][1][5] ^ A[3][2][5] ^ A[3][3][5] ^ A[3][4][5];
    assign C[3][6]     = A[3][0][6] ^ A[3][1][6] ^ A[3][2][6] ^ A[3][3][6] ^ A[3][4][6];
    assign C[3][7]     = A[3][0][7] ^ A[3][1][7] ^ A[3][2][7] ^ A[3][3][7] ^ A[3][4][7];
    assign C[3][8]     = A[3][0][8] ^ A[3][1][8] ^ A[3][2][8] ^ A[3][3][8] ^ A[3][4][8];
    assign C[3][9]     = A[3][0][9] ^ A[3][1][9] ^ A[3][2][9] ^ A[3][3][9] ^ A[3][4][9];
    assign C[3][10]     = A[3][0][10] ^ A[3][1][10] ^ A[3][2][10] ^ A[3][3][10] ^ A[3][4][10];
    assign C[3][11]     = A[3][0][11] ^ A[3][1][11] ^ A[3][2][11] ^ A[3][3][11] ^ A[3][4][11];
    assign C[3][12]     = A[3][0][12] ^ A[3][1][12] ^ A[3][2][12] ^ A[3][3][12] ^ A[3][4][12];
    assign C[3][13]     = A[3][0][13] ^ A[3][1][13] ^ A[3][2][13] ^ A[3][3][13] ^ A[3][4][13];
    assign C[3][14]     = A[3][0][14] ^ A[3][1][14] ^ A[3][2][14] ^ A[3][3][14] ^ A[3][4][14];
    assign C[3][15]     = A[3][0][15] ^ A[3][1][15] ^ A[3][2][15] ^ A[3][3][15] ^ A[3][4][15];
    assign C[3][16]     = A[3][0][16] ^ A[3][1][16] ^ A[3][2][16] ^ A[3][3][16] ^ A[3][4][16];
    assign C[3][17]     = A[3][0][17] ^ A[3][1][17] ^ A[3][2][17] ^ A[3][3][17] ^ A[3][4][17];
    assign C[3][18]     = A[3][0][18] ^ A[3][1][18] ^ A[3][2][18] ^ A[3][3][18] ^ A[3][4][18];
    assign C[3][19]     = A[3][0][19] ^ A[3][1][19] ^ A[3][2][19] ^ A[3][3][19] ^ A[3][4][19];
    assign C[3][20]     = A[3][0][20] ^ A[3][1][20] ^ A[3][2][20] ^ A[3][3][20] ^ A[3][4][20];
    assign C[3][21]     = A[3][0][21] ^ A[3][1][21] ^ A[3][2][21] ^ A[3][3][21] ^ A[3][4][21];
    assign C[3][22]     = A[3][0][22] ^ A[3][1][22] ^ A[3][2][22] ^ A[3][3][22] ^ A[3][4][22];
    assign C[3][23]     = A[3][0][23] ^ A[3][1][23] ^ A[3][2][23] ^ A[3][3][23] ^ A[3][4][23];
    assign C[3][24]     = A[3][0][24] ^ A[3][1][24] ^ A[3][2][24] ^ A[3][3][24] ^ A[3][4][24];
    assign C[3][25]     = A[3][0][25] ^ A[3][1][25] ^ A[3][2][25] ^ A[3][3][25] ^ A[3][4][25];
    assign C[3][26]     = A[3][0][26] ^ A[3][1][26] ^ A[3][2][26] ^ A[3][3][26] ^ A[3][4][26];
    assign C[3][27]     = A[3][0][27] ^ A[3][1][27] ^ A[3][2][27] ^ A[3][3][27] ^ A[3][4][27];
    assign C[3][28]     = A[3][0][28] ^ A[3][1][28] ^ A[3][2][28] ^ A[3][3][28] ^ A[3][4][28];
    assign C[3][29]     = A[3][0][29] ^ A[3][1][29] ^ A[3][2][29] ^ A[3][3][29] ^ A[3][4][29];
    assign C[3][30]     = A[3][0][30] ^ A[3][1][30] ^ A[3][2][30] ^ A[3][3][30] ^ A[3][4][30];
    assign C[3][31]     = A[3][0][31] ^ A[3][1][31] ^ A[3][2][31] ^ A[3][3][31] ^ A[3][4][31];
    assign C[3][32]     = A[3][0][32] ^ A[3][1][32] ^ A[3][2][32] ^ A[3][3][32] ^ A[3][4][32];
    assign C[3][33]     = A[3][0][33] ^ A[3][1][33] ^ A[3][2][33] ^ A[3][3][33] ^ A[3][4][33];
    assign C[3][34]     = A[3][0][34] ^ A[3][1][34] ^ A[3][2][34] ^ A[3][3][34] ^ A[3][4][34];
    assign C[3][35]     = A[3][0][35] ^ A[3][1][35] ^ A[3][2][35] ^ A[3][3][35] ^ A[3][4][35];
    assign C[3][36]     = A[3][0][36] ^ A[3][1][36] ^ A[3][2][36] ^ A[3][3][36] ^ A[3][4][36];
    assign C[3][37]     = A[3][0][37] ^ A[3][1][37] ^ A[3][2][37] ^ A[3][3][37] ^ A[3][4][37];
    assign C[3][38]     = A[3][0][38] ^ A[3][1][38] ^ A[3][2][38] ^ A[3][3][38] ^ A[3][4][38];
    assign C[3][39]     = A[3][0][39] ^ A[3][1][39] ^ A[3][2][39] ^ A[3][3][39] ^ A[3][4][39];
    assign C[3][40]     = A[3][0][40] ^ A[3][1][40] ^ A[3][2][40] ^ A[3][3][40] ^ A[3][4][40];
    assign C[3][41]     = A[3][0][41] ^ A[3][1][41] ^ A[3][2][41] ^ A[3][3][41] ^ A[3][4][41];
    assign C[3][42]     = A[3][0][42] ^ A[3][1][42] ^ A[3][2][42] ^ A[3][3][42] ^ A[3][4][42];
    assign C[3][43]     = A[3][0][43] ^ A[3][1][43] ^ A[3][2][43] ^ A[3][3][43] ^ A[3][4][43];
    assign C[3][44]     = A[3][0][44] ^ A[3][1][44] ^ A[3][2][44] ^ A[3][3][44] ^ A[3][4][44];
    assign C[3][45]     = A[3][0][45] ^ A[3][1][45] ^ A[3][2][45] ^ A[3][3][45] ^ A[3][4][45];
    assign C[3][46]     = A[3][0][46] ^ A[3][1][46] ^ A[3][2][46] ^ A[3][3][46] ^ A[3][4][46];
    assign C[3][47]     = A[3][0][47] ^ A[3][1][47] ^ A[3][2][47] ^ A[3][3][47] ^ A[3][4][47];
    assign C[3][48]     = A[3][0][48] ^ A[3][1][48] ^ A[3][2][48] ^ A[3][3][48] ^ A[3][4][48];
    assign C[3][49]     = A[3][0][49] ^ A[3][1][49] ^ A[3][2][49] ^ A[3][3][49] ^ A[3][4][49];
    assign C[3][50]     = A[3][0][50] ^ A[3][1][50] ^ A[3][2][50] ^ A[3][3][50] ^ A[3][4][50];
    assign C[3][51]     = A[3][0][51] ^ A[3][1][51] ^ A[3][2][51] ^ A[3][3][51] ^ A[3][4][51];
    assign C[3][52]     = A[3][0][52] ^ A[3][1][52] ^ A[3][2][52] ^ A[3][3][52] ^ A[3][4][52];
    assign C[3][53]     = A[3][0][53] ^ A[3][1][53] ^ A[3][2][53] ^ A[3][3][53] ^ A[3][4][53];
    assign C[3][54]     = A[3][0][54] ^ A[3][1][54] ^ A[3][2][54] ^ A[3][3][54] ^ A[3][4][54];
    assign C[3][55]     = A[3][0][55] ^ A[3][1][55] ^ A[3][2][55] ^ A[3][3][55] ^ A[3][4][55];
    assign C[3][56]     = A[3][0][56] ^ A[3][1][56] ^ A[3][2][56] ^ A[3][3][56] ^ A[3][4][56];
    assign C[3][57]     = A[3][0][57] ^ A[3][1][57] ^ A[3][2][57] ^ A[3][3][57] ^ A[3][4][57];
    assign C[3][58]     = A[3][0][58] ^ A[3][1][58] ^ A[3][2][58] ^ A[3][3][58] ^ A[3][4][58];
    assign C[3][59]     = A[3][0][59] ^ A[3][1][59] ^ A[3][2][59] ^ A[3][3][59] ^ A[3][4][59];
    assign C[3][60]     = A[3][0][60] ^ A[3][1][60] ^ A[3][2][60] ^ A[3][3][60] ^ A[3][4][60];
    assign C[3][61]     = A[3][0][61] ^ A[3][1][61] ^ A[3][2][61] ^ A[3][3][61] ^ A[3][4][61];
    assign C[3][62]     = A[3][0][62] ^ A[3][1][62] ^ A[3][2][62] ^ A[3][3][62] ^ A[3][4][62];
    assign C[3][63]     = A[3][0][63] ^ A[3][1][63] ^ A[3][2][63] ^ A[3][3][63] ^ A[3][4][63];
    assign C[4][0]     = A[4][0][0] ^ A[4][1][0] ^ A[4][2][0] ^ A[4][3][0] ^ A[4][4][0];
    assign C[4][1]     = A[4][0][1] ^ A[4][1][1] ^ A[4][2][1] ^ A[4][3][1] ^ A[4][4][1];
    assign C[4][2]     = A[4][0][2] ^ A[4][1][2] ^ A[4][2][2] ^ A[4][3][2] ^ A[4][4][2];
    assign C[4][3]     = A[4][0][3] ^ A[4][1][3] ^ A[4][2][3] ^ A[4][3][3] ^ A[4][4][3];
    assign C[4][4]     = A[4][0][4] ^ A[4][1][4] ^ A[4][2][4] ^ A[4][3][4] ^ A[4][4][4];
    assign C[4][5]     = A[4][0][5] ^ A[4][1][5] ^ A[4][2][5] ^ A[4][3][5] ^ A[4][4][5];
    assign C[4][6]     = A[4][0][6] ^ A[4][1][6] ^ A[4][2][6] ^ A[4][3][6] ^ A[4][4][6];
    assign C[4][7]     = A[4][0][7] ^ A[4][1][7] ^ A[4][2][7] ^ A[4][3][7] ^ A[4][4][7];
    assign C[4][8]     = A[4][0][8] ^ A[4][1][8] ^ A[4][2][8] ^ A[4][3][8] ^ A[4][4][8];
    assign C[4][9]     = A[4][0][9] ^ A[4][1][9] ^ A[4][2][9] ^ A[4][3][9] ^ A[4][4][9];
    assign C[4][10]     = A[4][0][10] ^ A[4][1][10] ^ A[4][2][10] ^ A[4][3][10] ^ A[4][4][10];
    assign C[4][11]     = A[4][0][11] ^ A[4][1][11] ^ A[4][2][11] ^ A[4][3][11] ^ A[4][4][11];
    assign C[4][12]     = A[4][0][12] ^ A[4][1][12] ^ A[4][2][12] ^ A[4][3][12] ^ A[4][4][12];
    assign C[4][13]     = A[4][0][13] ^ A[4][1][13] ^ A[4][2][13] ^ A[4][3][13] ^ A[4][4][13];
    assign C[4][14]     = A[4][0][14] ^ A[4][1][14] ^ A[4][2][14] ^ A[4][3][14] ^ A[4][4][14];
    assign C[4][15]     = A[4][0][15] ^ A[4][1][15] ^ A[4][2][15] ^ A[4][3][15] ^ A[4][4][15];
    assign C[4][16]     = A[4][0][16] ^ A[4][1][16] ^ A[4][2][16] ^ A[4][3][16] ^ A[4][4][16];
    assign C[4][17]     = A[4][0][17] ^ A[4][1][17] ^ A[4][2][17] ^ A[4][3][17] ^ A[4][4][17];
    assign C[4][18]     = A[4][0][18] ^ A[4][1][18] ^ A[4][2][18] ^ A[4][3][18] ^ A[4][4][18];
    assign C[4][19]     = A[4][0][19] ^ A[4][1][19] ^ A[4][2][19] ^ A[4][3][19] ^ A[4][4][19];
    assign C[4][20]     = A[4][0][20] ^ A[4][1][20] ^ A[4][2][20] ^ A[4][3][20] ^ A[4][4][20];
    assign C[4][21]     = A[4][0][21] ^ A[4][1][21] ^ A[4][2][21] ^ A[4][3][21] ^ A[4][4][21];
    assign C[4][22]     = A[4][0][22] ^ A[4][1][22] ^ A[4][2][22] ^ A[4][3][22] ^ A[4][4][22];
    assign C[4][23]     = A[4][0][23] ^ A[4][1][23] ^ A[4][2][23] ^ A[4][3][23] ^ A[4][4][23];
    assign C[4][24]     = A[4][0][24] ^ A[4][1][24] ^ A[4][2][24] ^ A[4][3][24] ^ A[4][4][24];
    assign C[4][25]     = A[4][0][25] ^ A[4][1][25] ^ A[4][2][25] ^ A[4][3][25] ^ A[4][4][25];
    assign C[4][26]     = A[4][0][26] ^ A[4][1][26] ^ A[4][2][26] ^ A[4][3][26] ^ A[4][4][26];
    assign C[4][27]     = A[4][0][27] ^ A[4][1][27] ^ A[4][2][27] ^ A[4][3][27] ^ A[4][4][27];
    assign C[4][28]     = A[4][0][28] ^ A[4][1][28] ^ A[4][2][28] ^ A[4][3][28] ^ A[4][4][28];
    assign C[4][29]     = A[4][0][29] ^ A[4][1][29] ^ A[4][2][29] ^ A[4][3][29] ^ A[4][4][29];
    assign C[4][30]     = A[4][0][30] ^ A[4][1][30] ^ A[4][2][30] ^ A[4][3][30] ^ A[4][4][30];
    assign C[4][31]     = A[4][0][31] ^ A[4][1][31] ^ A[4][2][31] ^ A[4][3][31] ^ A[4][4][31];
    assign C[4][32]     = A[4][0][32] ^ A[4][1][32] ^ A[4][2][32] ^ A[4][3][32] ^ A[4][4][32];
    assign C[4][33]     = A[4][0][33] ^ A[4][1][33] ^ A[4][2][33] ^ A[4][3][33] ^ A[4][4][33];
    assign C[4][34]     = A[4][0][34] ^ A[4][1][34] ^ A[4][2][34] ^ A[4][3][34] ^ A[4][4][34];
    assign C[4][35]     = A[4][0][35] ^ A[4][1][35] ^ A[4][2][35] ^ A[4][3][35] ^ A[4][4][35];
    assign C[4][36]     = A[4][0][36] ^ A[4][1][36] ^ A[4][2][36] ^ A[4][3][36] ^ A[4][4][36];
    assign C[4][37]     = A[4][0][37] ^ A[4][1][37] ^ A[4][2][37] ^ A[4][3][37] ^ A[4][4][37];
    assign C[4][38]     = A[4][0][38] ^ A[4][1][38] ^ A[4][2][38] ^ A[4][3][38] ^ A[4][4][38];
    assign C[4][39]     = A[4][0][39] ^ A[4][1][39] ^ A[4][2][39] ^ A[4][3][39] ^ A[4][4][39];
    assign C[4][40]     = A[4][0][40] ^ A[4][1][40] ^ A[4][2][40] ^ A[4][3][40] ^ A[4][4][40];
    assign C[4][41]     = A[4][0][41] ^ A[4][1][41] ^ A[4][2][41] ^ A[4][3][41] ^ A[4][4][41];
    assign C[4][42]     = A[4][0][42] ^ A[4][1][42] ^ A[4][2][42] ^ A[4][3][42] ^ A[4][4][42];
    assign C[4][43]     = A[4][0][43] ^ A[4][1][43] ^ A[4][2][43] ^ A[4][3][43] ^ A[4][4][43];
    assign C[4][44]     = A[4][0][44] ^ A[4][1][44] ^ A[4][2][44] ^ A[4][3][44] ^ A[4][4][44];
    assign C[4][45]     = A[4][0][45] ^ A[4][1][45] ^ A[4][2][45] ^ A[4][3][45] ^ A[4][4][45];
    assign C[4][46]     = A[4][0][46] ^ A[4][1][46] ^ A[4][2][46] ^ A[4][3][46] ^ A[4][4][46];
    assign C[4][47]     = A[4][0][47] ^ A[4][1][47] ^ A[4][2][47] ^ A[4][3][47] ^ A[4][4][47];
    assign C[4][48]     = A[4][0][48] ^ A[4][1][48] ^ A[4][2][48] ^ A[4][3][48] ^ A[4][4][48];
    assign C[4][49]     = A[4][0][49] ^ A[4][1][49] ^ A[4][2][49] ^ A[4][3][49] ^ A[4][4][49];
    assign C[4][50]     = A[4][0][50] ^ A[4][1][50] ^ A[4][2][50] ^ A[4][3][50] ^ A[4][4][50];
    assign C[4][51]     = A[4][0][51] ^ A[4][1][51] ^ A[4][2][51] ^ A[4][3][51] ^ A[4][4][51];
    assign C[4][52]     = A[4][0][52] ^ A[4][1][52] ^ A[4][2][52] ^ A[4][3][52] ^ A[4][4][52];
    assign C[4][53]     = A[4][0][53] ^ A[4][1][53] ^ A[4][2][53] ^ A[4][3][53] ^ A[4][4][53];
    assign C[4][54]     = A[4][0][54] ^ A[4][1][54] ^ A[4][2][54] ^ A[4][3][54] ^ A[4][4][54];
    assign C[4][55]     = A[4][0][55] ^ A[4][1][55] ^ A[4][2][55] ^ A[4][3][55] ^ A[4][4][55];
    assign C[4][56]     = A[4][0][56] ^ A[4][1][56] ^ A[4][2][56] ^ A[4][3][56] ^ A[4][4][56];
    assign C[4][57]     = A[4][0][57] ^ A[4][1][57] ^ A[4][2][57] ^ A[4][3][57] ^ A[4][4][57];
    assign C[4][58]     = A[4][0][58] ^ A[4][1][58] ^ A[4][2][58] ^ A[4][3][58] ^ A[4][4][58];
    assign C[4][59]     = A[4][0][59] ^ A[4][1][59] ^ A[4][2][59] ^ A[4][3][59] ^ A[4][4][59];
    assign C[4][60]     = A[4][0][60] ^ A[4][1][60] ^ A[4][2][60] ^ A[4][3][60] ^ A[4][4][60];
    assign C[4][61]     = A[4][0][61] ^ A[4][1][61] ^ A[4][2][61] ^ A[4][3][61] ^ A[4][4][61];
    assign C[4][62]     = A[4][0][62] ^ A[4][1][62] ^ A[4][2][62] ^ A[4][3][62] ^ A[4][4][62];
    assign C[4][63]     = A[4][0][63] ^ A[4][1][63] ^ A[4][2][63] ^ A[4][3][63] ^ A[4][4][63];

    // Step 2: Compute D[x][z]
    assign D[0][0]     = C[4][0] ^ C[1][63];
    assign D[0][1]     = C[4][1] ^ C[1][0];
    assign D[0][2]     = C[4][2] ^ C[1][1];
    assign D[0][3]     = C[4][3] ^ C[1][2];
    assign D[0][4]     = C[4][4] ^ C[1][3];
    assign D[0][5]     = C[4][5] ^ C[1][4];
    assign D[0][6]     = C[4][6] ^ C[1][5];
    assign D[0][7]     = C[4][7] ^ C[1][6];
    assign D[0][8]     = C[4][8] ^ C[1][7];
    assign D[0][9]     = C[4][9] ^ C[1][8];
    assign D[0][10]     = C[4][10] ^ C[1][9];
    assign D[0][11]     = C[4][11] ^ C[1][10];
    assign D[0][12]     = C[4][12] ^ C[1][11];
    assign D[0][13]     = C[4][13] ^ C[1][12];
    assign D[0][14]     = C[4][14] ^ C[1][13];
    assign D[0][15]     = C[4][15] ^ C[1][14];
    assign D[0][16]     = C[4][16] ^ C[1][15];
    assign D[0][17]     = C[4][17] ^ C[1][16];
    assign D[0][18]     = C[4][18] ^ C[1][17];
    assign D[0][19]     = C[4][19] ^ C[1][18];
    assign D[0][20]     = C[4][20] ^ C[1][19];
    assign D[0][21]     = C[4][21] ^ C[1][20];
    assign D[0][22]     = C[4][22] ^ C[1][21];
    assign D[0][23]     = C[4][23] ^ C[1][22];
    assign D[0][24]     = C[4][24] ^ C[1][23];
    assign D[0][25]     = C[4][25] ^ C[1][24];
    assign D[0][26]     = C[4][26] ^ C[1][25];
    assign D[0][27]     = C[4][27] ^ C[1][26];
    assign D[0][28]     = C[4][28] ^ C[1][27];
    assign D[0][29]     = C[4][29] ^ C[1][28];
    assign D[0][30]     = C[4][30] ^ C[1][29];
    assign D[0][31]     = C[4][31] ^ C[1][30];
    assign D[0][32]     = C[4][32] ^ C[1][31];
    assign D[0][33]     = C[4][33] ^ C[1][32];
    assign D[0][34]     = C[4][34] ^ C[1][33];
    assign D[0][35]     = C[4][35] ^ C[1][34];
    assign D[0][36]     = C[4][36] ^ C[1][35];
    assign D[0][37]     = C[4][37] ^ C[1][36];
    assign D[0][38]     = C[4][38] ^ C[1][37];
    assign D[0][39]     = C[4][39] ^ C[1][38];
    assign D[0][40]     = C[4][40] ^ C[1][39];
    assign D[0][41]     = C[4][41] ^ C[1][40];
    assign D[0][42]     = C[4][42] ^ C[1][41];
    assign D[0][43]     = C[4][43] ^ C[1][42];
    assign D[0][44]     = C[4][44] ^ C[1][43];
    assign D[0][45]     = C[4][45] ^ C[1][44];
    assign D[0][46]     = C[4][46] ^ C[1][45];
    assign D[0][47]     = C[4][47] ^ C[1][46];
    assign D[0][48]     = C[4][48] ^ C[1][47];
    assign D[0][49]     = C[4][49] ^ C[1][48];
    assign D[0][50]     = C[4][50] ^ C[1][49];
    assign D[0][51]     = C[4][51] ^ C[1][50];
    assign D[0][52]     = C[4][52] ^ C[1][51];
    assign D[0][53]     = C[4][53] ^ C[1][52];
    assign D[0][54]     = C[4][54] ^ C[1][53];
    assign D[0][55]     = C[4][55] ^ C[1][54];
    assign D[0][56]     = C[4][56] ^ C[1][55];
    assign D[0][57]     = C[4][57] ^ C[1][56];
    assign D[0][58]     = C[4][58] ^ C[1][57];
    assign D[0][59]     = C[4][59] ^ C[1][58];
    assign D[0][60]     = C[4][60] ^ C[1][59];
    assign D[0][61]     = C[4][61] ^ C[1][60];
    assign D[0][62]     = C[4][62] ^ C[1][61];
    assign D[0][63]     = C[4][63] ^ C[1][62];
    assign D[1][0]     = C[0][0] ^ C[2][63];
    assign D[1][1]     = C[0][1] ^ C[2][0];
    assign D[1][2]     = C[0][2] ^ C[2][1];
    assign D[1][3]     = C[0][3] ^ C[2][2];
    assign D[1][4]     = C[0][4] ^ C[2][3];
    assign D[1][5]     = C[0][5] ^ C[2][4];
    assign D[1][6]     = C[0][6] ^ C[2][5];
    assign D[1][7]     = C[0][7] ^ C[2][6];
    assign D[1][8]     = C[0][8] ^ C[2][7];
    assign D[1][9]     = C[0][9] ^ C[2][8];
    assign D[1][10]     = C[0][10] ^ C[2][9];
    assign D[1][11]     = C[0][11] ^ C[2][10];
    assign D[1][12]     = C[0][12] ^ C[2][11];
    assign D[1][13]     = C[0][13] ^ C[2][12];
    assign D[1][14]     = C[0][14] ^ C[2][13];
    assign D[1][15]     = C[0][15] ^ C[2][14];
    assign D[1][16]     = C[0][16] ^ C[2][15];
    assign D[1][17]     = C[0][17] ^ C[2][16];
    assign D[1][18]     = C[0][18] ^ C[2][17];
    assign D[1][19]     = C[0][19] ^ C[2][18];
    assign D[1][20]     = C[0][20] ^ C[2][19];
    assign D[1][21]     = C[0][21] ^ C[2][20];
    assign D[1][22]     = C[0][22] ^ C[2][21];
    assign D[1][23]     = C[0][23] ^ C[2][22];
    assign D[1][24]     = C[0][24] ^ C[2][23];
    assign D[1][25]     = C[0][25] ^ C[2][24];
    assign D[1][26]     = C[0][26] ^ C[2][25];
    assign D[1][27]     = C[0][27] ^ C[2][26];
    assign D[1][28]     = C[0][28] ^ C[2][27];
    assign D[1][29]     = C[0][29] ^ C[2][28];
    assign D[1][30]     = C[0][30] ^ C[2][29];
    assign D[1][31]     = C[0][31] ^ C[2][30];
    assign D[1][32]     = C[0][32] ^ C[2][31];
    assign D[1][33]     = C[0][33] ^ C[2][32];
    assign D[1][34]     = C[0][34] ^ C[2][33];
    assign D[1][35]     = C[0][35] ^ C[2][34];
    assign D[1][36]     = C[0][36] ^ C[2][35];
    assign D[1][37]     = C[0][37] ^ C[2][36];
    assign D[1][38]     = C[0][38] ^ C[2][37];
    assign D[1][39]     = C[0][39] ^ C[2][38];
    assign D[1][40]     = C[0][40] ^ C[2][39];
    assign D[1][41]     = C[0][41] ^ C[2][40];
    assign D[1][42]     = C[0][42] ^ C[2][41];
    assign D[1][43]     = C[0][43] ^ C[2][42];
    assign D[1][44]     = C[0][44] ^ C[2][43];
    assign D[1][45]     = C[0][45] ^ C[2][44];
    assign D[1][46]     = C[0][46] ^ C[2][45];
    assign D[1][47]     = C[0][47] ^ C[2][46];
    assign D[1][48]     = C[0][48] ^ C[2][47];
    assign D[1][49]     = C[0][49] ^ C[2][48];
    assign D[1][50]     = C[0][50] ^ C[2][49];
    assign D[1][51]     = C[0][51] ^ C[2][50];
    assign D[1][52]     = C[0][52] ^ C[2][51];
    assign D[1][53]     = C[0][53] ^ C[2][52];
    assign D[1][54]     = C[0][54] ^ C[2][53];
    assign D[1][55]     = C[0][55] ^ C[2][54];
    assign D[1][56]     = C[0][56] ^ C[2][55];
    assign D[1][57]     = C[0][57] ^ C[2][56];
    assign D[1][58]     = C[0][58] ^ C[2][57];
    assign D[1][59]     = C[0][59] ^ C[2][58];
    assign D[1][60]     = C[0][60] ^ C[2][59];
    assign D[1][61]     = C[0][61] ^ C[2][60];
    assign D[1][62]     = C[0][62] ^ C[2][61];
    assign D[1][63]     = C[0][63] ^ C[2][62];
    assign D[2][0]     = C[1][0] ^ C[3][63];
    assign D[2][1]     = C[1][1] ^ C[3][0];
    assign D[2][2]     = C[1][2] ^ C[3][1];
    assign D[2][3]     = C[1][3] ^ C[3][2];
    assign D[2][4]     = C[1][4] ^ C[3][3];
    assign D[2][5]     = C[1][5] ^ C[3][4];
    assign D[2][6]     = C[1][6] ^ C[3][5];
    assign D[2][7]     = C[1][7] ^ C[3][6];
    assign D[2][8]     = C[1][8] ^ C[3][7];
    assign D[2][9]     = C[1][9] ^ C[3][8];
    assign D[2][10]     = C[1][10] ^ C[3][9];
    assign D[2][11]     = C[1][11] ^ C[3][10];
    assign D[2][12]     = C[1][12] ^ C[3][11];
    assign D[2][13]     = C[1][13] ^ C[3][12];
    assign D[2][14]     = C[1][14] ^ C[3][13];
    assign D[2][15]     = C[1][15] ^ C[3][14];
    assign D[2][16]     = C[1][16] ^ C[3][15];
    assign D[2][17]     = C[1][17] ^ C[3][16];
    assign D[2][18]     = C[1][18] ^ C[3][17];
    assign D[2][19]     = C[1][19] ^ C[3][18];
    assign D[2][20]     = C[1][20] ^ C[3][19];
    assign D[2][21]     = C[1][21] ^ C[3][20];
    assign D[2][22]     = C[1][22] ^ C[3][21];
    assign D[2][23]     = C[1][23] ^ C[3][22];
    assign D[2][24]     = C[1][24] ^ C[3][23];
    assign D[2][25]     = C[1][25] ^ C[3][24];
    assign D[2][26]     = C[1][26] ^ C[3][25];
    assign D[2][27]     = C[1][27] ^ C[3][26];
    assign D[2][28]     = C[1][28] ^ C[3][27];
    assign D[2][29]     = C[1][29] ^ C[3][28];
    assign D[2][30]     = C[1][30] ^ C[3][29];
    assign D[2][31]     = C[1][31] ^ C[3][30];
    assign D[2][32]     = C[1][32] ^ C[3][31];
    assign D[2][33]     = C[1][33] ^ C[3][32];
    assign D[2][34]     = C[1][34] ^ C[3][33];
    assign D[2][35]     = C[1][35] ^ C[3][34];
    assign D[2][36]     = C[1][36] ^ C[3][35];
    assign D[2][37]     = C[1][37] ^ C[3][36];
    assign D[2][38]     = C[1][38] ^ C[3][37];
    assign D[2][39]     = C[1][39] ^ C[3][38];
    assign D[2][40]     = C[1][40] ^ C[3][39];
    assign D[2][41]     = C[1][41] ^ C[3][40];
    assign D[2][42]     = C[1][42] ^ C[3][41];
    assign D[2][43]     = C[1][43] ^ C[3][42];
    assign D[2][44]     = C[1][44] ^ C[3][43];
    assign D[2][45]     = C[1][45] ^ C[3][44];
    assign D[2][46]     = C[1][46] ^ C[3][45];
    assign D[2][47]     = C[1][47] ^ C[3][46];
    assign D[2][48]     = C[1][48] ^ C[3][47];
    assign D[2][49]     = C[1][49] ^ C[3][48];
    assign D[2][50]     = C[1][50] ^ C[3][49];
    assign D[2][51]     = C[1][51] ^ C[3][50];
    assign D[2][52]     = C[1][52] ^ C[3][51];
    assign D[2][53]     = C[1][53] ^ C[3][52];
    assign D[2][54]     = C[1][54] ^ C[3][53];
    assign D[2][55]     = C[1][55] ^ C[3][54];
    assign D[2][56]     = C[1][56] ^ C[3][55];
    assign D[2][57]     = C[1][57] ^ C[3][56];
    assign D[2][58]     = C[1][58] ^ C[3][57];
    assign D[2][59]     = C[1][59] ^ C[3][58];
    assign D[2][60]     = C[1][60] ^ C[3][59];
    assign D[2][61]     = C[1][61] ^ C[3][60];
    assign D[2][62]     = C[1][62] ^ C[3][61];
    assign D[2][63]     = C[1][63] ^ C[3][62];
    assign D[3][0]     = C[2][0] ^ C[4][63];
    assign D[3][1]     = C[2][1] ^ C[4][0];
    assign D[3][2]     = C[2][2] ^ C[4][1];
    assign D[3][3]     = C[2][3] ^ C[4][2];
    assign D[3][4]     = C[2][4] ^ C[4][3];
    assign D[3][5]     = C[2][5] ^ C[4][4];
    assign D[3][6]     = C[2][6] ^ C[4][5];
    assign D[3][7]     = C[2][7] ^ C[4][6];
    assign D[3][8]     = C[2][8] ^ C[4][7];
    assign D[3][9]     = C[2][9] ^ C[4][8];
    assign D[3][10]     = C[2][10] ^ C[4][9];
    assign D[3][11]     = C[2][11] ^ C[4][10];
    assign D[3][12]     = C[2][12] ^ C[4][11];
    assign D[3][13]     = C[2][13] ^ C[4][12];
    assign D[3][14]     = C[2][14] ^ C[4][13];
    assign D[3][15]     = C[2][15] ^ C[4][14];
    assign D[3][16]     = C[2][16] ^ C[4][15];
    assign D[3][17]     = C[2][17] ^ C[4][16];
    assign D[3][18]     = C[2][18] ^ C[4][17];
    assign D[3][19]     = C[2][19] ^ C[4][18];
    assign D[3][20]     = C[2][20] ^ C[4][19];
    assign D[3][21]     = C[2][21] ^ C[4][20];
    assign D[3][22]     = C[2][22] ^ C[4][21];
    assign D[3][23]     = C[2][23] ^ C[4][22];
    assign D[3][24]     = C[2][24] ^ C[4][23];
    assign D[3][25]     = C[2][25] ^ C[4][24];
    assign D[3][26]     = C[2][26] ^ C[4][25];
    assign D[3][27]     = C[2][27] ^ C[4][26];
    assign D[3][28]     = C[2][28] ^ C[4][27];
    assign D[3][29]     = C[2][29] ^ C[4][28];
    assign D[3][30]     = C[2][30] ^ C[4][29];
    assign D[3][31]     = C[2][31] ^ C[4][30];
    assign D[3][32]     = C[2][32] ^ C[4][31];
    assign D[3][33]     = C[2][33] ^ C[4][32];
    assign D[3][34]     = C[2][34] ^ C[4][33];
    assign D[3][35]     = C[2][35] ^ C[4][34];
    assign D[3][36]     = C[2][36] ^ C[4][35];
    assign D[3][37]     = C[2][37] ^ C[4][36];
    assign D[3][38]     = C[2][38] ^ C[4][37];
    assign D[3][39]     = C[2][39] ^ C[4][38];
    assign D[3][40]     = C[2][40] ^ C[4][39];
    assign D[3][41]     = C[2][41] ^ C[4][40];
    assign D[3][42]     = C[2][42] ^ C[4][41];
    assign D[3][43]     = C[2][43] ^ C[4][42];
    assign D[3][44]     = C[2][44] ^ C[4][43];
    assign D[3][45]     = C[2][45] ^ C[4][44];
    assign D[3][46]     = C[2][46] ^ C[4][45];
    assign D[3][47]     = C[2][47] ^ C[4][46];
    assign D[3][48]     = C[2][48] ^ C[4][47];
    assign D[3][49]     = C[2][49] ^ C[4][48];
    assign D[3][50]     = C[2][50] ^ C[4][49];
    assign D[3][51]     = C[2][51] ^ C[4][50];
    assign D[3][52]     = C[2][52] ^ C[4][51];
    assign D[3][53]     = C[2][53] ^ C[4][52];
    assign D[3][54]     = C[2][54] ^ C[4][53];
    assign D[3][55]     = C[2][55] ^ C[4][54];
    assign D[3][56]     = C[2][56] ^ C[4][55];
    assign D[3][57]     = C[2][57] ^ C[4][56];
    assign D[3][58]     = C[2][58] ^ C[4][57];
    assign D[3][59]     = C[2][59] ^ C[4][58];
    assign D[3][60]     = C[2][60] ^ C[4][59];
    assign D[3][61]     = C[2][61] ^ C[4][60];
    assign D[3][62]     = C[2][62] ^ C[4][61];
    assign D[3][63]     = C[2][63] ^ C[4][62];
    assign D[4][0]     = C[3][0] ^ C[0][63];
    assign D[4][1]     = C[3][1] ^ C[0][0];
    assign D[4][2]     = C[3][2] ^ C[0][1];
    assign D[4][3]     = C[3][3] ^ C[0][2];
    assign D[4][4]     = C[3][4] ^ C[0][3];
    assign D[4][5]     = C[3][5] ^ C[0][4];
    assign D[4][6]     = C[3][6] ^ C[0][5];
    assign D[4][7]     = C[3][7] ^ C[0][6];
    assign D[4][8]     = C[3][8] ^ C[0][7];
    assign D[4][9]     = C[3][9] ^ C[0][8];
    assign D[4][10]     = C[3][10] ^ C[0][9];
    assign D[4][11]     = C[3][11] ^ C[0][10];
    assign D[4][12]     = C[3][12] ^ C[0][11];
    assign D[4][13]     = C[3][13] ^ C[0][12];
    assign D[4][14]     = C[3][14] ^ C[0][13];
    assign D[4][15]     = C[3][15] ^ C[0][14];
    assign D[4][16]     = C[3][16] ^ C[0][15];
    assign D[4][17]     = C[3][17] ^ C[0][16];
    assign D[4][18]     = C[3][18] ^ C[0][17];
    assign D[4][19]     = C[3][19] ^ C[0][18];
    assign D[4][20]     = C[3][20] ^ C[0][19];
    assign D[4][21]     = C[3][21] ^ C[0][20];
    assign D[4][22]     = C[3][22] ^ C[0][21];
    assign D[4][23]     = C[3][23] ^ C[0][22];
    assign D[4][24]     = C[3][24] ^ C[0][23];
    assign D[4][25]     = C[3][25] ^ C[0][24];
    assign D[4][26]     = C[3][26] ^ C[0][25];
    assign D[4][27]     = C[3][27] ^ C[0][26];
    assign D[4][28]     = C[3][28] ^ C[0][27];
    assign D[4][29]     = C[3][29] ^ C[0][28];
    assign D[4][30]     = C[3][30] ^ C[0][29];
    assign D[4][31]     = C[3][31] ^ C[0][30];
    assign D[4][32]     = C[3][32] ^ C[0][31];
    assign D[4][33]     = C[3][33] ^ C[0][32];
    assign D[4][34]     = C[3][34] ^ C[0][33];
    assign D[4][35]     = C[3][35] ^ C[0][34];
    assign D[4][36]     = C[3][36] ^ C[0][35];
    assign D[4][37]     = C[3][37] ^ C[0][36];
    assign D[4][38]     = C[3][38] ^ C[0][37];
    assign D[4][39]     = C[3][39] ^ C[0][38];
    assign D[4][40]     = C[3][40] ^ C[0][39];
    assign D[4][41]     = C[3][41] ^ C[0][40];
    assign D[4][42]     = C[3][42] ^ C[0][41];
    assign D[4][43]     = C[3][43] ^ C[0][42];
    assign D[4][44]     = C[3][44] ^ C[0][43];
    assign D[4][45]     = C[3][45] ^ C[0][44];
    assign D[4][46]     = C[3][46] ^ C[0][45];
    assign D[4][47]     = C[3][47] ^ C[0][46];
    assign D[4][48]     = C[3][48] ^ C[0][47];
    assign D[4][49]     = C[3][49] ^ C[0][48];
    assign D[4][50]     = C[3][50] ^ C[0][49];
    assign D[4][51]     = C[3][51] ^ C[0][50];
    assign D[4][52]     = C[3][52] ^ C[0][51];
    assign D[4][53]     = C[3][53] ^ C[0][52];
    assign D[4][54]     = C[3][54] ^ C[0][53];
    assign D[4][55]     = C[3][55] ^ C[0][54];
    assign D[4][56]     = C[3][56] ^ C[0][55];
    assign D[4][57]     = C[3][57] ^ C[0][56];
    assign D[4][58]     = C[3][58] ^ C[0][57];
    assign D[4][59]     = C[3][59] ^ C[0][58];
    assign D[4][60]     = C[3][60] ^ C[0][59];
    assign D[4][61]     = C[3][61] ^ C[0][60];
    assign D[4][62]     = C[3][62] ^ C[0][61];
    assign D[4][63]     = C[3][63] ^ C[0][62];

    // Step 3: Compute A_theta[x][y][z] = A[x][y][z] ^ D[x][z]
    assign A_theta[0][0][0]  = A[0][0][0] ^ D[0][0];
    assign A_theta[0][0][1]  = A[0][0][1] ^ D[0][1];
    assign A_theta[0][0][2]  = A[0][0][2] ^ D[0][2];
    assign A_theta[0][0][3]  = A[0][0][3] ^ D[0][3];
    assign A_theta[0][0][4]  = A[0][0][4] ^ D[0][4];
    assign A_theta[0][0][5]  = A[0][0][5] ^ D[0][5];
    assign A_theta[0][0][6]  = A[0][0][6] ^ D[0][6];
    assign A_theta[0][0][7]  = A[0][0][7] ^ D[0][7];
    assign A_theta[0][0][8]  = A[0][0][8] ^ D[0][8];
    assign A_theta[0][0][9]  = A[0][0][9] ^ D[0][9];
    assign A_theta[0][0][10]  = A[0][0][10] ^ D[0][10];
    assign A_theta[0][0][11]  = A[0][0][11] ^ D[0][11];
    assign A_theta[0][0][12]  = A[0][0][12] ^ D[0][12];
    assign A_theta[0][0][13]  = A[0][0][13] ^ D[0][13];
    assign A_theta[0][0][14]  = A[0][0][14] ^ D[0][14];
    assign A_theta[0][0][15]  = A[0][0][15] ^ D[0][15];
    assign A_theta[0][0][16]  = A[0][0][16] ^ D[0][16];
    assign A_theta[0][0][17]  = A[0][0][17] ^ D[0][17];
    assign A_theta[0][0][18]  = A[0][0][18] ^ D[0][18];
    assign A_theta[0][0][19]  = A[0][0][19] ^ D[0][19];
    assign A_theta[0][0][20]  = A[0][0][20] ^ D[0][20];
    assign A_theta[0][0][21]  = A[0][0][21] ^ D[0][21];
    assign A_theta[0][0][22]  = A[0][0][22] ^ D[0][22];
    assign A_theta[0][0][23]  = A[0][0][23] ^ D[0][23];
    assign A_theta[0][0][24]  = A[0][0][24] ^ D[0][24];
    assign A_theta[0][0][25]  = A[0][0][25] ^ D[0][25];
    assign A_theta[0][0][26]  = A[0][0][26] ^ D[0][26];
    assign A_theta[0][0][27]  = A[0][0][27] ^ D[0][27];
    assign A_theta[0][0][28]  = A[0][0][28] ^ D[0][28];
    assign A_theta[0][0][29]  = A[0][0][29] ^ D[0][29];
    assign A_theta[0][0][30]  = A[0][0][30] ^ D[0][30];
    assign A_theta[0][0][31]  = A[0][0][31] ^ D[0][31];
    assign A_theta[0][0][32]  = A[0][0][32] ^ D[0][32];
    assign A_theta[0][0][33]  = A[0][0][33] ^ D[0][33];
    assign A_theta[0][0][34]  = A[0][0][34] ^ D[0][34];
    assign A_theta[0][0][35]  = A[0][0][35] ^ D[0][35];
    assign A_theta[0][0][36]  = A[0][0][36] ^ D[0][36];
    assign A_theta[0][0][37]  = A[0][0][37] ^ D[0][37];
    assign A_theta[0][0][38]  = A[0][0][38] ^ D[0][38];
    assign A_theta[0][0][39]  = A[0][0][39] ^ D[0][39];
    assign A_theta[0][0][40]  = A[0][0][40] ^ D[0][40];
    assign A_theta[0][0][41]  = A[0][0][41] ^ D[0][41];
    assign A_theta[0][0][42]  = A[0][0][42] ^ D[0][42];
    assign A_theta[0][0][43]  = A[0][0][43] ^ D[0][43];
    assign A_theta[0][0][44]  = A[0][0][44] ^ D[0][44];
    assign A_theta[0][0][45]  = A[0][0][45] ^ D[0][45];
    assign A_theta[0][0][46]  = A[0][0][46] ^ D[0][46];
    assign A_theta[0][0][47]  = A[0][0][47] ^ D[0][47];
    assign A_theta[0][0][48]  = A[0][0][48] ^ D[0][48];
    assign A_theta[0][0][49]  = A[0][0][49] ^ D[0][49];
    assign A_theta[0][0][50]  = A[0][0][50] ^ D[0][50];
    assign A_theta[0][0][51]  = A[0][0][51] ^ D[0][51];
    assign A_theta[0][0][52]  = A[0][0][52] ^ D[0][52];
    assign A_theta[0][0][53]  = A[0][0][53] ^ D[0][53];
    assign A_theta[0][0][54]  = A[0][0][54] ^ D[0][54];
    assign A_theta[0][0][55]  = A[0][0][55] ^ D[0][55];
    assign A_theta[0][0][56]  = A[0][0][56] ^ D[0][56];
    assign A_theta[0][0][57]  = A[0][0][57] ^ D[0][57];
    assign A_theta[0][0][58]  = A[0][0][58] ^ D[0][58];
    assign A_theta[0][0][59]  = A[0][0][59] ^ D[0][59];
    assign A_theta[0][0][60]  = A[0][0][60] ^ D[0][60];
    assign A_theta[0][0][61]  = A[0][0][61] ^ D[0][61];
    assign A_theta[0][0][62]  = A[0][0][62] ^ D[0][62];
    assign A_theta[0][0][63]  = A[0][0][63] ^ D[0][63];
    assign A_theta[0][1][0]  = A[0][1][0] ^ D[0][0];
    assign A_theta[0][1][1]  = A[0][1][1] ^ D[0][1];
    assign A_theta[0][1][2]  = A[0][1][2] ^ D[0][2];
    assign A_theta[0][1][3]  = A[0][1][3] ^ D[0][3];
    assign A_theta[0][1][4]  = A[0][1][4] ^ D[0][4];
    assign A_theta[0][1][5]  = A[0][1][5] ^ D[0][5];
    assign A_theta[0][1][6]  = A[0][1][6] ^ D[0][6];
    assign A_theta[0][1][7]  = A[0][1][7] ^ D[0][7];
    assign A_theta[0][1][8]  = A[0][1][8] ^ D[0][8];
    assign A_theta[0][1][9]  = A[0][1][9] ^ D[0][9];
    assign A_theta[0][1][10]  = A[0][1][10] ^ D[0][10];
    assign A_theta[0][1][11]  = A[0][1][11] ^ D[0][11];
    assign A_theta[0][1][12]  = A[0][1][12] ^ D[0][12];
    assign A_theta[0][1][13]  = A[0][1][13] ^ D[0][13];
    assign A_theta[0][1][14]  = A[0][1][14] ^ D[0][14];
    assign A_theta[0][1][15]  = A[0][1][15] ^ D[0][15];
    assign A_theta[0][1][16]  = A[0][1][16] ^ D[0][16];
    assign A_theta[0][1][17]  = A[0][1][17] ^ D[0][17];
    assign A_theta[0][1][18]  = A[0][1][18] ^ D[0][18];
    assign A_theta[0][1][19]  = A[0][1][19] ^ D[0][19];
    assign A_theta[0][1][20]  = A[0][1][20] ^ D[0][20];
    assign A_theta[0][1][21]  = A[0][1][21] ^ D[0][21];
    assign A_theta[0][1][22]  = A[0][1][22] ^ D[0][22];
    assign A_theta[0][1][23]  = A[0][1][23] ^ D[0][23];
    assign A_theta[0][1][24]  = A[0][1][24] ^ D[0][24];
    assign A_theta[0][1][25]  = A[0][1][25] ^ D[0][25];
    assign A_theta[0][1][26]  = A[0][1][26] ^ D[0][26];
    assign A_theta[0][1][27]  = A[0][1][27] ^ D[0][27];
    assign A_theta[0][1][28]  = A[0][1][28] ^ D[0][28];
    assign A_theta[0][1][29]  = A[0][1][29] ^ D[0][29];
    assign A_theta[0][1][30]  = A[0][1][30] ^ D[0][30];
    assign A_theta[0][1][31]  = A[0][1][31] ^ D[0][31];
    assign A_theta[0][1][32]  = A[0][1][32] ^ D[0][32];
    assign A_theta[0][1][33]  = A[0][1][33] ^ D[0][33];
    assign A_theta[0][1][34]  = A[0][1][34] ^ D[0][34];
    assign A_theta[0][1][35]  = A[0][1][35] ^ D[0][35];
    assign A_theta[0][1][36]  = A[0][1][36] ^ D[0][36];
    assign A_theta[0][1][37]  = A[0][1][37] ^ D[0][37];
    assign A_theta[0][1][38]  = A[0][1][38] ^ D[0][38];
    assign A_theta[0][1][39]  = A[0][1][39] ^ D[0][39];
    assign A_theta[0][1][40]  = A[0][1][40] ^ D[0][40];
    assign A_theta[0][1][41]  = A[0][1][41] ^ D[0][41];
    assign A_theta[0][1][42]  = A[0][1][42] ^ D[0][42];
    assign A_theta[0][1][43]  = A[0][1][43] ^ D[0][43];
    assign A_theta[0][1][44]  = A[0][1][44] ^ D[0][44];
    assign A_theta[0][1][45]  = A[0][1][45] ^ D[0][45];
    assign A_theta[0][1][46]  = A[0][1][46] ^ D[0][46];
    assign A_theta[0][1][47]  = A[0][1][47] ^ D[0][47];
    assign A_theta[0][1][48]  = A[0][1][48] ^ D[0][48];
    assign A_theta[0][1][49]  = A[0][1][49] ^ D[0][49];
    assign A_theta[0][1][50]  = A[0][1][50] ^ D[0][50];
    assign A_theta[0][1][51]  = A[0][1][51] ^ D[0][51];
    assign A_theta[0][1][52]  = A[0][1][52] ^ D[0][52];
    assign A_theta[0][1][53]  = A[0][1][53] ^ D[0][53];
    assign A_theta[0][1][54]  = A[0][1][54] ^ D[0][54];
    assign A_theta[0][1][55]  = A[0][1][55] ^ D[0][55];
    assign A_theta[0][1][56]  = A[0][1][56] ^ D[0][56];
    assign A_theta[0][1][57]  = A[0][1][57] ^ D[0][57];
    assign A_theta[0][1][58]  = A[0][1][58] ^ D[0][58];
    assign A_theta[0][1][59]  = A[0][1][59] ^ D[0][59];
    assign A_theta[0][1][60]  = A[0][1][60] ^ D[0][60];
    assign A_theta[0][1][61]  = A[0][1][61] ^ D[0][61];
    assign A_theta[0][1][62]  = A[0][1][62] ^ D[0][62];
    assign A_theta[0][1][63]  = A[0][1][63] ^ D[0][63];
    assign A_theta[0][2][0]  = A[0][2][0] ^ D[0][0];
    assign A_theta[0][2][1]  = A[0][2][1] ^ D[0][1];
    assign A_theta[0][2][2]  = A[0][2][2] ^ D[0][2];
    assign A_theta[0][2][3]  = A[0][2][3] ^ D[0][3];
    assign A_theta[0][2][4]  = A[0][2][4] ^ D[0][4];
    assign A_theta[0][2][5]  = A[0][2][5] ^ D[0][5];
    assign A_theta[0][2][6]  = A[0][2][6] ^ D[0][6];
    assign A_theta[0][2][7]  = A[0][2][7] ^ D[0][7];
    assign A_theta[0][2][8]  = A[0][2][8] ^ D[0][8];
    assign A_theta[0][2][9]  = A[0][2][9] ^ D[0][9];
    assign A_theta[0][2][10]  = A[0][2][10] ^ D[0][10];
    assign A_theta[0][2][11]  = A[0][2][11] ^ D[0][11];
    assign A_theta[0][2][12]  = A[0][2][12] ^ D[0][12];
    assign A_theta[0][2][13]  = A[0][2][13] ^ D[0][13];
    assign A_theta[0][2][14]  = A[0][2][14] ^ D[0][14];
    assign A_theta[0][2][15]  = A[0][2][15] ^ D[0][15];
    assign A_theta[0][2][16]  = A[0][2][16] ^ D[0][16];
    assign A_theta[0][2][17]  = A[0][2][17] ^ D[0][17];
    assign A_theta[0][2][18]  = A[0][2][18] ^ D[0][18];
    assign A_theta[0][2][19]  = A[0][2][19] ^ D[0][19];
    assign A_theta[0][2][20]  = A[0][2][20] ^ D[0][20];
    assign A_theta[0][2][21]  = A[0][2][21] ^ D[0][21];
    assign A_theta[0][2][22]  = A[0][2][22] ^ D[0][22];
    assign A_theta[0][2][23]  = A[0][2][23] ^ D[0][23];
    assign A_theta[0][2][24]  = A[0][2][24] ^ D[0][24];
    assign A_theta[0][2][25]  = A[0][2][25] ^ D[0][25];
    assign A_theta[0][2][26]  = A[0][2][26] ^ D[0][26];
    assign A_theta[0][2][27]  = A[0][2][27] ^ D[0][27];
    assign A_theta[0][2][28]  = A[0][2][28] ^ D[0][28];
    assign A_theta[0][2][29]  = A[0][2][29] ^ D[0][29];
    assign A_theta[0][2][30]  = A[0][2][30] ^ D[0][30];
    assign A_theta[0][2][31]  = A[0][2][31] ^ D[0][31];
    assign A_theta[0][2][32]  = A[0][2][32] ^ D[0][32];
    assign A_theta[0][2][33]  = A[0][2][33] ^ D[0][33];
    assign A_theta[0][2][34]  = A[0][2][34] ^ D[0][34];
    assign A_theta[0][2][35]  = A[0][2][35] ^ D[0][35];
    assign A_theta[0][2][36]  = A[0][2][36] ^ D[0][36];
    assign A_theta[0][2][37]  = A[0][2][37] ^ D[0][37];
    assign A_theta[0][2][38]  = A[0][2][38] ^ D[0][38];
    assign A_theta[0][2][39]  = A[0][2][39] ^ D[0][39];
    assign A_theta[0][2][40]  = A[0][2][40] ^ D[0][40];
    assign A_theta[0][2][41]  = A[0][2][41] ^ D[0][41];
    assign A_theta[0][2][42]  = A[0][2][42] ^ D[0][42];
    assign A_theta[0][2][43]  = A[0][2][43] ^ D[0][43];
    assign A_theta[0][2][44]  = A[0][2][44] ^ D[0][44];
    assign A_theta[0][2][45]  = A[0][2][45] ^ D[0][45];
    assign A_theta[0][2][46]  = A[0][2][46] ^ D[0][46];
    assign A_theta[0][2][47]  = A[0][2][47] ^ D[0][47];
    assign A_theta[0][2][48]  = A[0][2][48] ^ D[0][48];
    assign A_theta[0][2][49]  = A[0][2][49] ^ D[0][49];
    assign A_theta[0][2][50]  = A[0][2][50] ^ D[0][50];
    assign A_theta[0][2][51]  = A[0][2][51] ^ D[0][51];
    assign A_theta[0][2][52]  = A[0][2][52] ^ D[0][52];
    assign A_theta[0][2][53]  = A[0][2][53] ^ D[0][53];
    assign A_theta[0][2][54]  = A[0][2][54] ^ D[0][54];
    assign A_theta[0][2][55]  = A[0][2][55] ^ D[0][55];
    assign A_theta[0][2][56]  = A[0][2][56] ^ D[0][56];
    assign A_theta[0][2][57]  = A[0][2][57] ^ D[0][57];
    assign A_theta[0][2][58]  = A[0][2][58] ^ D[0][58];
    assign A_theta[0][2][59]  = A[0][2][59] ^ D[0][59];
    assign A_theta[0][2][60]  = A[0][2][60] ^ D[0][60];
    assign A_theta[0][2][61]  = A[0][2][61] ^ D[0][61];
    assign A_theta[0][2][62]  = A[0][2][62] ^ D[0][62];
    assign A_theta[0][2][63]  = A[0][2][63] ^ D[0][63];
    assign A_theta[0][3][0]  = A[0][3][0] ^ D[0][0];
    assign A_theta[0][3][1]  = A[0][3][1] ^ D[0][1];
    assign A_theta[0][3][2]  = A[0][3][2] ^ D[0][2];
    assign A_theta[0][3][3]  = A[0][3][3] ^ D[0][3];
    assign A_theta[0][3][4]  = A[0][3][4] ^ D[0][4];
    assign A_theta[0][3][5]  = A[0][3][5] ^ D[0][5];
    assign A_theta[0][3][6]  = A[0][3][6] ^ D[0][6];
    assign A_theta[0][3][7]  = A[0][3][7] ^ D[0][7];
    assign A_theta[0][3][8]  = A[0][3][8] ^ D[0][8];
    assign A_theta[0][3][9]  = A[0][3][9] ^ D[0][9];
    assign A_theta[0][3][10]  = A[0][3][10] ^ D[0][10];
    assign A_theta[0][3][11]  = A[0][3][11] ^ D[0][11];
    assign A_theta[0][3][12]  = A[0][3][12] ^ D[0][12];
    assign A_theta[0][3][13]  = A[0][3][13] ^ D[0][13];
    assign A_theta[0][3][14]  = A[0][3][14] ^ D[0][14];
    assign A_theta[0][3][15]  = A[0][3][15] ^ D[0][15];
    assign A_theta[0][3][16]  = A[0][3][16] ^ D[0][16];
    assign A_theta[0][3][17]  = A[0][3][17] ^ D[0][17];
    assign A_theta[0][3][18]  = A[0][3][18] ^ D[0][18];
    assign A_theta[0][3][19]  = A[0][3][19] ^ D[0][19];
    assign A_theta[0][3][20]  = A[0][3][20] ^ D[0][20];
    assign A_theta[0][3][21]  = A[0][3][21] ^ D[0][21];
    assign A_theta[0][3][22]  = A[0][3][22] ^ D[0][22];
    assign A_theta[0][3][23]  = A[0][3][23] ^ D[0][23];
    assign A_theta[0][3][24]  = A[0][3][24] ^ D[0][24];
    assign A_theta[0][3][25]  = A[0][3][25] ^ D[0][25];
    assign A_theta[0][3][26]  = A[0][3][26] ^ D[0][26];
    assign A_theta[0][3][27]  = A[0][3][27] ^ D[0][27];
    assign A_theta[0][3][28]  = A[0][3][28] ^ D[0][28];
    assign A_theta[0][3][29]  = A[0][3][29] ^ D[0][29];
    assign A_theta[0][3][30]  = A[0][3][30] ^ D[0][30];
    assign A_theta[0][3][31]  = A[0][3][31] ^ D[0][31];
    assign A_theta[0][3][32]  = A[0][3][32] ^ D[0][32];
    assign A_theta[0][3][33]  = A[0][3][33] ^ D[0][33];
    assign A_theta[0][3][34]  = A[0][3][34] ^ D[0][34];
    assign A_theta[0][3][35]  = A[0][3][35] ^ D[0][35];
    assign A_theta[0][3][36]  = A[0][3][36] ^ D[0][36];
    assign A_theta[0][3][37]  = A[0][3][37] ^ D[0][37];
    assign A_theta[0][3][38]  = A[0][3][38] ^ D[0][38];
    assign A_theta[0][3][39]  = A[0][3][39] ^ D[0][39];
    assign A_theta[0][3][40]  = A[0][3][40] ^ D[0][40];
    assign A_theta[0][3][41]  = A[0][3][41] ^ D[0][41];
    assign A_theta[0][3][42]  = A[0][3][42] ^ D[0][42];
    assign A_theta[0][3][43]  = A[0][3][43] ^ D[0][43];
    assign A_theta[0][3][44]  = A[0][3][44] ^ D[0][44];
    assign A_theta[0][3][45]  = A[0][3][45] ^ D[0][45];
    assign A_theta[0][3][46]  = A[0][3][46] ^ D[0][46];
    assign A_theta[0][3][47]  = A[0][3][47] ^ D[0][47];
    assign A_theta[0][3][48]  = A[0][3][48] ^ D[0][48];
    assign A_theta[0][3][49]  = A[0][3][49] ^ D[0][49];
    assign A_theta[0][3][50]  = A[0][3][50] ^ D[0][50];
    assign A_theta[0][3][51]  = A[0][3][51] ^ D[0][51];
    assign A_theta[0][3][52]  = A[0][3][52] ^ D[0][52];
    assign A_theta[0][3][53]  = A[0][3][53] ^ D[0][53];
    assign A_theta[0][3][54]  = A[0][3][54] ^ D[0][54];
    assign A_theta[0][3][55]  = A[0][3][55] ^ D[0][55];
    assign A_theta[0][3][56]  = A[0][3][56] ^ D[0][56];
    assign A_theta[0][3][57]  = A[0][3][57] ^ D[0][57];
    assign A_theta[0][3][58]  = A[0][3][58] ^ D[0][58];
    assign A_theta[0][3][59]  = A[0][3][59] ^ D[0][59];
    assign A_theta[0][3][60]  = A[0][3][60] ^ D[0][60];
    assign A_theta[0][3][61]  = A[0][3][61] ^ D[0][61];
    assign A_theta[0][3][62]  = A[0][3][62] ^ D[0][62];
    assign A_theta[0][3][63]  = A[0][3][63] ^ D[0][63];
    assign A_theta[0][4][0]  = A[0][4][0] ^ D[0][0];
    assign A_theta[0][4][1]  = A[0][4][1] ^ D[0][1];
    assign A_theta[0][4][2]  = A[0][4][2] ^ D[0][2];
    assign A_theta[0][4][3]  = A[0][4][3] ^ D[0][3];
    assign A_theta[0][4][4]  = A[0][4][4] ^ D[0][4];
    assign A_theta[0][4][5]  = A[0][4][5] ^ D[0][5];
    assign A_theta[0][4][6]  = A[0][4][6] ^ D[0][6];
    assign A_theta[0][4][7]  = A[0][4][7] ^ D[0][7];
    assign A_theta[0][4][8]  = A[0][4][8] ^ D[0][8];
    assign A_theta[0][4][9]  = A[0][4][9] ^ D[0][9];
    assign A_theta[0][4][10]  = A[0][4][10] ^ D[0][10];
    assign A_theta[0][4][11]  = A[0][4][11] ^ D[0][11];
    assign A_theta[0][4][12]  = A[0][4][12] ^ D[0][12];
    assign A_theta[0][4][13]  = A[0][4][13] ^ D[0][13];
    assign A_theta[0][4][14]  = A[0][4][14] ^ D[0][14];
    assign A_theta[0][4][15]  = A[0][4][15] ^ D[0][15];
    assign A_theta[0][4][16]  = A[0][4][16] ^ D[0][16];
    assign A_theta[0][4][17]  = A[0][4][17] ^ D[0][17];
    assign A_theta[0][4][18]  = A[0][4][18] ^ D[0][18];
    assign A_theta[0][4][19]  = A[0][4][19] ^ D[0][19];
    assign A_theta[0][4][20]  = A[0][4][20] ^ D[0][20];
    assign A_theta[0][4][21]  = A[0][4][21] ^ D[0][21];
    assign A_theta[0][4][22]  = A[0][4][22] ^ D[0][22];
    assign A_theta[0][4][23]  = A[0][4][23] ^ D[0][23];
    assign A_theta[0][4][24]  = A[0][4][24] ^ D[0][24];
    assign A_theta[0][4][25]  = A[0][4][25] ^ D[0][25];
    assign A_theta[0][4][26]  = A[0][4][26] ^ D[0][26];
    assign A_theta[0][4][27]  = A[0][4][27] ^ D[0][27];
    assign A_theta[0][4][28]  = A[0][4][28] ^ D[0][28];
    assign A_theta[0][4][29]  = A[0][4][29] ^ D[0][29];
    assign A_theta[0][4][30]  = A[0][4][30] ^ D[0][30];
    assign A_theta[0][4][31]  = A[0][4][31] ^ D[0][31];
    assign A_theta[0][4][32]  = A[0][4][32] ^ D[0][32];
    assign A_theta[0][4][33]  = A[0][4][33] ^ D[0][33];
    assign A_theta[0][4][34]  = A[0][4][34] ^ D[0][34];
    assign A_theta[0][4][35]  = A[0][4][35] ^ D[0][35];
    assign A_theta[0][4][36]  = A[0][4][36] ^ D[0][36];
    assign A_theta[0][4][37]  = A[0][4][37] ^ D[0][37];
    assign A_theta[0][4][38]  = A[0][4][38] ^ D[0][38];
    assign A_theta[0][4][39]  = A[0][4][39] ^ D[0][39];
    assign A_theta[0][4][40]  = A[0][4][40] ^ D[0][40];
    assign A_theta[0][4][41]  = A[0][4][41] ^ D[0][41];
    assign A_theta[0][4][42]  = A[0][4][42] ^ D[0][42];
    assign A_theta[0][4][43]  = A[0][4][43] ^ D[0][43];
    assign A_theta[0][4][44]  = A[0][4][44] ^ D[0][44];
    assign A_theta[0][4][45]  = A[0][4][45] ^ D[0][45];
    assign A_theta[0][4][46]  = A[0][4][46] ^ D[0][46];
    assign A_theta[0][4][47]  = A[0][4][47] ^ D[0][47];
    assign A_theta[0][4][48]  = A[0][4][48] ^ D[0][48];
    assign A_theta[0][4][49]  = A[0][4][49] ^ D[0][49];
    assign A_theta[0][4][50]  = A[0][4][50] ^ D[0][50];
    assign A_theta[0][4][51]  = A[0][4][51] ^ D[0][51];
    assign A_theta[0][4][52]  = A[0][4][52] ^ D[0][52];
    assign A_theta[0][4][53]  = A[0][4][53] ^ D[0][53];
    assign A_theta[0][4][54]  = A[0][4][54] ^ D[0][54];
    assign A_theta[0][4][55]  = A[0][4][55] ^ D[0][55];
    assign A_theta[0][4][56]  = A[0][4][56] ^ D[0][56];
    assign A_theta[0][4][57]  = A[0][4][57] ^ D[0][57];
    assign A_theta[0][4][58]  = A[0][4][58] ^ D[0][58];
    assign A_theta[0][4][59]  = A[0][4][59] ^ D[0][59];
    assign A_theta[0][4][60]  = A[0][4][60] ^ D[0][60];
    assign A_theta[0][4][61]  = A[0][4][61] ^ D[0][61];
    assign A_theta[0][4][62]  = A[0][4][62] ^ D[0][62];
    assign A_theta[0][4][63]  = A[0][4][63] ^ D[0][63];
    assign A_theta[1][0][0]  = A[1][0][0] ^ D[1][0];
    assign A_theta[1][0][1]  = A[1][0][1] ^ D[1][1];
    assign A_theta[1][0][2]  = A[1][0][2] ^ D[1][2];
    assign A_theta[1][0][3]  = A[1][0][3] ^ D[1][3];
    assign A_theta[1][0][4]  = A[1][0][4] ^ D[1][4];
    assign A_theta[1][0][5]  = A[1][0][5] ^ D[1][5];
    assign A_theta[1][0][6]  = A[1][0][6] ^ D[1][6];
    assign A_theta[1][0][7]  = A[1][0][7] ^ D[1][7];
    assign A_theta[1][0][8]  = A[1][0][8] ^ D[1][8];
    assign A_theta[1][0][9]  = A[1][0][9] ^ D[1][9];
    assign A_theta[1][0][10]  = A[1][0][10] ^ D[1][10];
    assign A_theta[1][0][11]  = A[1][0][11] ^ D[1][11];
    assign A_theta[1][0][12]  = A[1][0][12] ^ D[1][12];
    assign A_theta[1][0][13]  = A[1][0][13] ^ D[1][13];
    assign A_theta[1][0][14]  = A[1][0][14] ^ D[1][14];
    assign A_theta[1][0][15]  = A[1][0][15] ^ D[1][15];
    assign A_theta[1][0][16]  = A[1][0][16] ^ D[1][16];
    assign A_theta[1][0][17]  = A[1][0][17] ^ D[1][17];
    assign A_theta[1][0][18]  = A[1][0][18] ^ D[1][18];
    assign A_theta[1][0][19]  = A[1][0][19] ^ D[1][19];
    assign A_theta[1][0][20]  = A[1][0][20] ^ D[1][20];
    assign A_theta[1][0][21]  = A[1][0][21] ^ D[1][21];
    assign A_theta[1][0][22]  = A[1][0][22] ^ D[1][22];
    assign A_theta[1][0][23]  = A[1][0][23] ^ D[1][23];
    assign A_theta[1][0][24]  = A[1][0][24] ^ D[1][24];
    assign A_theta[1][0][25]  = A[1][0][25] ^ D[1][25];
    assign A_theta[1][0][26]  = A[1][0][26] ^ D[1][26];
    assign A_theta[1][0][27]  = A[1][0][27] ^ D[1][27];
    assign A_theta[1][0][28]  = A[1][0][28] ^ D[1][28];
    assign A_theta[1][0][29]  = A[1][0][29] ^ D[1][29];
    assign A_theta[1][0][30]  = A[1][0][30] ^ D[1][30];
    assign A_theta[1][0][31]  = A[1][0][31] ^ D[1][31];
    assign A_theta[1][0][32]  = A[1][0][32] ^ D[1][32];
    assign A_theta[1][0][33]  = A[1][0][33] ^ D[1][33];
    assign A_theta[1][0][34]  = A[1][0][34] ^ D[1][34];
    assign A_theta[1][0][35]  = A[1][0][35] ^ D[1][35];
    assign A_theta[1][0][36]  = A[1][0][36] ^ D[1][36];
    assign A_theta[1][0][37]  = A[1][0][37] ^ D[1][37];
    assign A_theta[1][0][38]  = A[1][0][38] ^ D[1][38];
    assign A_theta[1][0][39]  = A[1][0][39] ^ D[1][39];
    assign A_theta[1][0][40]  = A[1][0][40] ^ D[1][40];
    assign A_theta[1][0][41]  = A[1][0][41] ^ D[1][41];
    assign A_theta[1][0][42]  = A[1][0][42] ^ D[1][42];
    assign A_theta[1][0][43]  = A[1][0][43] ^ D[1][43];
    assign A_theta[1][0][44]  = A[1][0][44] ^ D[1][44];
    assign A_theta[1][0][45]  = A[1][0][45] ^ D[1][45];
    assign A_theta[1][0][46]  = A[1][0][46] ^ D[1][46];
    assign A_theta[1][0][47]  = A[1][0][47] ^ D[1][47];
    assign A_theta[1][0][48]  = A[1][0][48] ^ D[1][48];
    assign A_theta[1][0][49]  = A[1][0][49] ^ D[1][49];
    assign A_theta[1][0][50]  = A[1][0][50] ^ D[1][50];
    assign A_theta[1][0][51]  = A[1][0][51] ^ D[1][51];
    assign A_theta[1][0][52]  = A[1][0][52] ^ D[1][52];
    assign A_theta[1][0][53]  = A[1][0][53] ^ D[1][53];
    assign A_theta[1][0][54]  = A[1][0][54] ^ D[1][54];
    assign A_theta[1][0][55]  = A[1][0][55] ^ D[1][55];
    assign A_theta[1][0][56]  = A[1][0][56] ^ D[1][56];
    assign A_theta[1][0][57]  = A[1][0][57] ^ D[1][57];
    assign A_theta[1][0][58]  = A[1][0][58] ^ D[1][58];
    assign A_theta[1][0][59]  = A[1][0][59] ^ D[1][59];
    assign A_theta[1][0][60]  = A[1][0][60] ^ D[1][60];
    assign A_theta[1][0][61]  = A[1][0][61] ^ D[1][61];
    assign A_theta[1][0][62]  = A[1][0][62] ^ D[1][62];
    assign A_theta[1][0][63]  = A[1][0][63] ^ D[1][63];
    assign A_theta[1][1][0]  = A[1][1][0] ^ D[1][0];
    assign A_theta[1][1][1]  = A[1][1][1] ^ D[1][1];
    assign A_theta[1][1][2]  = A[1][1][2] ^ D[1][2];
    assign A_theta[1][1][3]  = A[1][1][3] ^ D[1][3];
    assign A_theta[1][1][4]  = A[1][1][4] ^ D[1][4];
    assign A_theta[1][1][5]  = A[1][1][5] ^ D[1][5];
    assign A_theta[1][1][6]  = A[1][1][6] ^ D[1][6];
    assign A_theta[1][1][7]  = A[1][1][7] ^ D[1][7];
    assign A_theta[1][1][8]  = A[1][1][8] ^ D[1][8];
    assign A_theta[1][1][9]  = A[1][1][9] ^ D[1][9];
    assign A_theta[1][1][10]  = A[1][1][10] ^ D[1][10];
    assign A_theta[1][1][11]  = A[1][1][11] ^ D[1][11];
    assign A_theta[1][1][12]  = A[1][1][12] ^ D[1][12];
    assign A_theta[1][1][13]  = A[1][1][13] ^ D[1][13];
    assign A_theta[1][1][14]  = A[1][1][14] ^ D[1][14];
    assign A_theta[1][1][15]  = A[1][1][15] ^ D[1][15];
    assign A_theta[1][1][16]  = A[1][1][16] ^ D[1][16];
    assign A_theta[1][1][17]  = A[1][1][17] ^ D[1][17];
    assign A_theta[1][1][18]  = A[1][1][18] ^ D[1][18];
    assign A_theta[1][1][19]  = A[1][1][19] ^ D[1][19];
    assign A_theta[1][1][20]  = A[1][1][20] ^ D[1][20];
    assign A_theta[1][1][21]  = A[1][1][21] ^ D[1][21];
    assign A_theta[1][1][22]  = A[1][1][22] ^ D[1][22];
    assign A_theta[1][1][23]  = A[1][1][23] ^ D[1][23];
    assign A_theta[1][1][24]  = A[1][1][24] ^ D[1][24];
    assign A_theta[1][1][25]  = A[1][1][25] ^ D[1][25];
    assign A_theta[1][1][26]  = A[1][1][26] ^ D[1][26];
    assign A_theta[1][1][27]  = A[1][1][27] ^ D[1][27];
    assign A_theta[1][1][28]  = A[1][1][28] ^ D[1][28];
    assign A_theta[1][1][29]  = A[1][1][29] ^ D[1][29];
    assign A_theta[1][1][30]  = A[1][1][30] ^ D[1][30];
    assign A_theta[1][1][31]  = A[1][1][31] ^ D[1][31];
    assign A_theta[1][1][32]  = A[1][1][32] ^ D[1][32];
    assign A_theta[1][1][33]  = A[1][1][33] ^ D[1][33];
    assign A_theta[1][1][34]  = A[1][1][34] ^ D[1][34];
    assign A_theta[1][1][35]  = A[1][1][35] ^ D[1][35];
    assign A_theta[1][1][36]  = A[1][1][36] ^ D[1][36];
    assign A_theta[1][1][37]  = A[1][1][37] ^ D[1][37];
    assign A_theta[1][1][38]  = A[1][1][38] ^ D[1][38];
    assign A_theta[1][1][39]  = A[1][1][39] ^ D[1][39];
    assign A_theta[1][1][40]  = A[1][1][40] ^ D[1][40];
    assign A_theta[1][1][41]  = A[1][1][41] ^ D[1][41];
    assign A_theta[1][1][42]  = A[1][1][42] ^ D[1][42];
    assign A_theta[1][1][43]  = A[1][1][43] ^ D[1][43];
    assign A_theta[1][1][44]  = A[1][1][44] ^ D[1][44];
    assign A_theta[1][1][45]  = A[1][1][45] ^ D[1][45];
    assign A_theta[1][1][46]  = A[1][1][46] ^ D[1][46];
    assign A_theta[1][1][47]  = A[1][1][47] ^ D[1][47];
    assign A_theta[1][1][48]  = A[1][1][48] ^ D[1][48];
    assign A_theta[1][1][49]  = A[1][1][49] ^ D[1][49];
    assign A_theta[1][1][50]  = A[1][1][50] ^ D[1][50];
    assign A_theta[1][1][51]  = A[1][1][51] ^ D[1][51];
    assign A_theta[1][1][52]  = A[1][1][52] ^ D[1][52];
    assign A_theta[1][1][53]  = A[1][1][53] ^ D[1][53];
    assign A_theta[1][1][54]  = A[1][1][54] ^ D[1][54];
    assign A_theta[1][1][55]  = A[1][1][55] ^ D[1][55];
    assign A_theta[1][1][56]  = A[1][1][56] ^ D[1][56];
    assign A_theta[1][1][57]  = A[1][1][57] ^ D[1][57];
    assign A_theta[1][1][58]  = A[1][1][58] ^ D[1][58];
    assign A_theta[1][1][59]  = A[1][1][59] ^ D[1][59];
    assign A_theta[1][1][60]  = A[1][1][60] ^ D[1][60];
    assign A_theta[1][1][61]  = A[1][1][61] ^ D[1][61];
    assign A_theta[1][1][62]  = A[1][1][62] ^ D[1][62];
    assign A_theta[1][1][63]  = A[1][1][63] ^ D[1][63];
    assign A_theta[1][2][0]  = A[1][2][0] ^ D[1][0];
    assign A_theta[1][2][1]  = A[1][2][1] ^ D[1][1];
    assign A_theta[1][2][2]  = A[1][2][2] ^ D[1][2];
    assign A_theta[1][2][3]  = A[1][2][3] ^ D[1][3];
    assign A_theta[1][2][4]  = A[1][2][4] ^ D[1][4];
    assign A_theta[1][2][5]  = A[1][2][5] ^ D[1][5];
    assign A_theta[1][2][6]  = A[1][2][6] ^ D[1][6];
    assign A_theta[1][2][7]  = A[1][2][7] ^ D[1][7];
    assign A_theta[1][2][8]  = A[1][2][8] ^ D[1][8];
    assign A_theta[1][2][9]  = A[1][2][9] ^ D[1][9];
    assign A_theta[1][2][10]  = A[1][2][10] ^ D[1][10];
    assign A_theta[1][2][11]  = A[1][2][11] ^ D[1][11];
    assign A_theta[1][2][12]  = A[1][2][12] ^ D[1][12];
    assign A_theta[1][2][13]  = A[1][2][13] ^ D[1][13];
    assign A_theta[1][2][14]  = A[1][2][14] ^ D[1][14];
    assign A_theta[1][2][15]  = A[1][2][15] ^ D[1][15];
    assign A_theta[1][2][16]  = A[1][2][16] ^ D[1][16];
    assign A_theta[1][2][17]  = A[1][2][17] ^ D[1][17];
    assign A_theta[1][2][18]  = A[1][2][18] ^ D[1][18];
    assign A_theta[1][2][19]  = A[1][2][19] ^ D[1][19];
    assign A_theta[1][2][20]  = A[1][2][20] ^ D[1][20];
    assign A_theta[1][2][21]  = A[1][2][21] ^ D[1][21];
    assign A_theta[1][2][22]  = A[1][2][22] ^ D[1][22];
    assign A_theta[1][2][23]  = A[1][2][23] ^ D[1][23];
    assign A_theta[1][2][24]  = A[1][2][24] ^ D[1][24];
    assign A_theta[1][2][25]  = A[1][2][25] ^ D[1][25];
    assign A_theta[1][2][26]  = A[1][2][26] ^ D[1][26];
    assign A_theta[1][2][27]  = A[1][2][27] ^ D[1][27];
    assign A_theta[1][2][28]  = A[1][2][28] ^ D[1][28];
    assign A_theta[1][2][29]  = A[1][2][29] ^ D[1][29];
    assign A_theta[1][2][30]  = A[1][2][30] ^ D[1][30];
    assign A_theta[1][2][31]  = A[1][2][31] ^ D[1][31];
    assign A_theta[1][2][32]  = A[1][2][32] ^ D[1][32];
    assign A_theta[1][2][33]  = A[1][2][33] ^ D[1][33];
    assign A_theta[1][2][34]  = A[1][2][34] ^ D[1][34];
    assign A_theta[1][2][35]  = A[1][2][35] ^ D[1][35];
    assign A_theta[1][2][36]  = A[1][2][36] ^ D[1][36];
    assign A_theta[1][2][37]  = A[1][2][37] ^ D[1][37];
    assign A_theta[1][2][38]  = A[1][2][38] ^ D[1][38];
    assign A_theta[1][2][39]  = A[1][2][39] ^ D[1][39];
    assign A_theta[1][2][40]  = A[1][2][40] ^ D[1][40];
    assign A_theta[1][2][41]  = A[1][2][41] ^ D[1][41];
    assign A_theta[1][2][42]  = A[1][2][42] ^ D[1][42];
    assign A_theta[1][2][43]  = A[1][2][43] ^ D[1][43];
    assign A_theta[1][2][44]  = A[1][2][44] ^ D[1][44];
    assign A_theta[1][2][45]  = A[1][2][45] ^ D[1][45];
    assign A_theta[1][2][46]  = A[1][2][46] ^ D[1][46];
    assign A_theta[1][2][47]  = A[1][2][47] ^ D[1][47];
    assign A_theta[1][2][48]  = A[1][2][48] ^ D[1][48];
    assign A_theta[1][2][49]  = A[1][2][49] ^ D[1][49];
    assign A_theta[1][2][50]  = A[1][2][50] ^ D[1][50];
    assign A_theta[1][2][51]  = A[1][2][51] ^ D[1][51];
    assign A_theta[1][2][52]  = A[1][2][52] ^ D[1][52];
    assign A_theta[1][2][53]  = A[1][2][53] ^ D[1][53];
    assign A_theta[1][2][54]  = A[1][2][54] ^ D[1][54];
    assign A_theta[1][2][55]  = A[1][2][55] ^ D[1][55];
    assign A_theta[1][2][56]  = A[1][2][56] ^ D[1][56];
    assign A_theta[1][2][57]  = A[1][2][57] ^ D[1][57];
    assign A_theta[1][2][58]  = A[1][2][58] ^ D[1][58];
    assign A_theta[1][2][59]  = A[1][2][59] ^ D[1][59];
    assign A_theta[1][2][60]  = A[1][2][60] ^ D[1][60];
    assign A_theta[1][2][61]  = A[1][2][61] ^ D[1][61];
    assign A_theta[1][2][62]  = A[1][2][62] ^ D[1][62];
    assign A_theta[1][2][63]  = A[1][2][63] ^ D[1][63];
    assign A_theta[1][3][0]  = A[1][3][0] ^ D[1][0];
    assign A_theta[1][3][1]  = A[1][3][1] ^ D[1][1];
    assign A_theta[1][3][2]  = A[1][3][2] ^ D[1][2];
    assign A_theta[1][3][3]  = A[1][3][3] ^ D[1][3];
    assign A_theta[1][3][4]  = A[1][3][4] ^ D[1][4];
    assign A_theta[1][3][5]  = A[1][3][5] ^ D[1][5];
    assign A_theta[1][3][6]  = A[1][3][6] ^ D[1][6];
    assign A_theta[1][3][7]  = A[1][3][7] ^ D[1][7];
    assign A_theta[1][3][8]  = A[1][3][8] ^ D[1][8];
    assign A_theta[1][3][9]  = A[1][3][9] ^ D[1][9];
    assign A_theta[1][3][10]  = A[1][3][10] ^ D[1][10];
    assign A_theta[1][3][11]  = A[1][3][11] ^ D[1][11];
    assign A_theta[1][3][12]  = A[1][3][12] ^ D[1][12];
    assign A_theta[1][3][13]  = A[1][3][13] ^ D[1][13];
    assign A_theta[1][3][14]  = A[1][3][14] ^ D[1][14];
    assign A_theta[1][3][15]  = A[1][3][15] ^ D[1][15];
    assign A_theta[1][3][16]  = A[1][3][16] ^ D[1][16];
    assign A_theta[1][3][17]  = A[1][3][17] ^ D[1][17];
    assign A_theta[1][3][18]  = A[1][3][18] ^ D[1][18];
    assign A_theta[1][3][19]  = A[1][3][19] ^ D[1][19];
    assign A_theta[1][3][20]  = A[1][3][20] ^ D[1][20];
    assign A_theta[1][3][21]  = A[1][3][21] ^ D[1][21];
    assign A_theta[1][3][22]  = A[1][3][22] ^ D[1][22];
    assign A_theta[1][3][23]  = A[1][3][23] ^ D[1][23];
    assign A_theta[1][3][24]  = A[1][3][24] ^ D[1][24];
    assign A_theta[1][3][25]  = A[1][3][25] ^ D[1][25];
    assign A_theta[1][3][26]  = A[1][3][26] ^ D[1][26];
    assign A_theta[1][3][27]  = A[1][3][27] ^ D[1][27];
    assign A_theta[1][3][28]  = A[1][3][28] ^ D[1][28];
    assign A_theta[1][3][29]  = A[1][3][29] ^ D[1][29];
    assign A_theta[1][3][30]  = A[1][3][30] ^ D[1][30];
    assign A_theta[1][3][31]  = A[1][3][31] ^ D[1][31];
    assign A_theta[1][3][32]  = A[1][3][32] ^ D[1][32];
    assign A_theta[1][3][33]  = A[1][3][33] ^ D[1][33];
    assign A_theta[1][3][34]  = A[1][3][34] ^ D[1][34];
    assign A_theta[1][3][35]  = A[1][3][35] ^ D[1][35];
    assign A_theta[1][3][36]  = A[1][3][36] ^ D[1][36];
    assign A_theta[1][3][37]  = A[1][3][37] ^ D[1][37];
    assign A_theta[1][3][38]  = A[1][3][38] ^ D[1][38];
    assign A_theta[1][3][39]  = A[1][3][39] ^ D[1][39];
    assign A_theta[1][3][40]  = A[1][3][40] ^ D[1][40];
    assign A_theta[1][3][41]  = A[1][3][41] ^ D[1][41];
    assign A_theta[1][3][42]  = A[1][3][42] ^ D[1][42];
    assign A_theta[1][3][43]  = A[1][3][43] ^ D[1][43];
    assign A_theta[1][3][44]  = A[1][3][44] ^ D[1][44];
    assign A_theta[1][3][45]  = A[1][3][45] ^ D[1][45];
    assign A_theta[1][3][46]  = A[1][3][46] ^ D[1][46];
    assign A_theta[1][3][47]  = A[1][3][47] ^ D[1][47];
    assign A_theta[1][3][48]  = A[1][3][48] ^ D[1][48];
    assign A_theta[1][3][49]  = A[1][3][49] ^ D[1][49];
    assign A_theta[1][3][50]  = A[1][3][50] ^ D[1][50];
    assign A_theta[1][3][51]  = A[1][3][51] ^ D[1][51];
    assign A_theta[1][3][52]  = A[1][3][52] ^ D[1][52];
    assign A_theta[1][3][53]  = A[1][3][53] ^ D[1][53];
    assign A_theta[1][3][54]  = A[1][3][54] ^ D[1][54];
    assign A_theta[1][3][55]  = A[1][3][55] ^ D[1][55];
    assign A_theta[1][3][56]  = A[1][3][56] ^ D[1][56];
    assign A_theta[1][3][57]  = A[1][3][57] ^ D[1][57];
    assign A_theta[1][3][58]  = A[1][3][58] ^ D[1][58];
    assign A_theta[1][3][59]  = A[1][3][59] ^ D[1][59];
    assign A_theta[1][3][60]  = A[1][3][60] ^ D[1][60];
    assign A_theta[1][3][61]  = A[1][3][61] ^ D[1][61];
    assign A_theta[1][3][62]  = A[1][3][62] ^ D[1][62];
    assign A_theta[1][3][63]  = A[1][3][63] ^ D[1][63];
    assign A_theta[1][4][0]  = A[1][4][0] ^ D[1][0];
    assign A_theta[1][4][1]  = A[1][4][1] ^ D[1][1];
    assign A_theta[1][4][2]  = A[1][4][2] ^ D[1][2];
    assign A_theta[1][4][3]  = A[1][4][3] ^ D[1][3];
    assign A_theta[1][4][4]  = A[1][4][4] ^ D[1][4];
    assign A_theta[1][4][5]  = A[1][4][5] ^ D[1][5];
    assign A_theta[1][4][6]  = A[1][4][6] ^ D[1][6];
    assign A_theta[1][4][7]  = A[1][4][7] ^ D[1][7];
    assign A_theta[1][4][8]  = A[1][4][8] ^ D[1][8];
    assign A_theta[1][4][9]  = A[1][4][9] ^ D[1][9];
    assign A_theta[1][4][10]  = A[1][4][10] ^ D[1][10];
    assign A_theta[1][4][11]  = A[1][4][11] ^ D[1][11];
    assign A_theta[1][4][12]  = A[1][4][12] ^ D[1][12];
    assign A_theta[1][4][13]  = A[1][4][13] ^ D[1][13];
    assign A_theta[1][4][14]  = A[1][4][14] ^ D[1][14];
    assign A_theta[1][4][15]  = A[1][4][15] ^ D[1][15];
    assign A_theta[1][4][16]  = A[1][4][16] ^ D[1][16];
    assign A_theta[1][4][17]  = A[1][4][17] ^ D[1][17];
    assign A_theta[1][4][18]  = A[1][4][18] ^ D[1][18];
    assign A_theta[1][4][19]  = A[1][4][19] ^ D[1][19];
    assign A_theta[1][4][20]  = A[1][4][20] ^ D[1][20];
    assign A_theta[1][4][21]  = A[1][4][21] ^ D[1][21];
    assign A_theta[1][4][22]  = A[1][4][22] ^ D[1][22];
    assign A_theta[1][4][23]  = A[1][4][23] ^ D[1][23];
    assign A_theta[1][4][24]  = A[1][4][24] ^ D[1][24];
    assign A_theta[1][4][25]  = A[1][4][25] ^ D[1][25];
    assign A_theta[1][4][26]  = A[1][4][26] ^ D[1][26];
    assign A_theta[1][4][27]  = A[1][4][27] ^ D[1][27];
    assign A_theta[1][4][28]  = A[1][4][28] ^ D[1][28];
    assign A_theta[1][4][29]  = A[1][4][29] ^ D[1][29];
    assign A_theta[1][4][30]  = A[1][4][30] ^ D[1][30];
    assign A_theta[1][4][31]  = A[1][4][31] ^ D[1][31];
    assign A_theta[1][4][32]  = A[1][4][32] ^ D[1][32];
    assign A_theta[1][4][33]  = A[1][4][33] ^ D[1][33];
    assign A_theta[1][4][34]  = A[1][4][34] ^ D[1][34];
    assign A_theta[1][4][35]  = A[1][4][35] ^ D[1][35];
    assign A_theta[1][4][36]  = A[1][4][36] ^ D[1][36];
    assign A_theta[1][4][37]  = A[1][4][37] ^ D[1][37];
    assign A_theta[1][4][38]  = A[1][4][38] ^ D[1][38];
    assign A_theta[1][4][39]  = A[1][4][39] ^ D[1][39];
    assign A_theta[1][4][40]  = A[1][4][40] ^ D[1][40];
    assign A_theta[1][4][41]  = A[1][4][41] ^ D[1][41];
    assign A_theta[1][4][42]  = A[1][4][42] ^ D[1][42];
    assign A_theta[1][4][43]  = A[1][4][43] ^ D[1][43];
    assign A_theta[1][4][44]  = A[1][4][44] ^ D[1][44];
    assign A_theta[1][4][45]  = A[1][4][45] ^ D[1][45];
    assign A_theta[1][4][46]  = A[1][4][46] ^ D[1][46];
    assign A_theta[1][4][47]  = A[1][4][47] ^ D[1][47];
    assign A_theta[1][4][48]  = A[1][4][48] ^ D[1][48];
    assign A_theta[1][4][49]  = A[1][4][49] ^ D[1][49];
    assign A_theta[1][4][50]  = A[1][4][50] ^ D[1][50];
    assign A_theta[1][4][51]  = A[1][4][51] ^ D[1][51];
    assign A_theta[1][4][52]  = A[1][4][52] ^ D[1][52];
    assign A_theta[1][4][53]  = A[1][4][53] ^ D[1][53];
    assign A_theta[1][4][54]  = A[1][4][54] ^ D[1][54];
    assign A_theta[1][4][55]  = A[1][4][55] ^ D[1][55];
    assign A_theta[1][4][56]  = A[1][4][56] ^ D[1][56];
    assign A_theta[1][4][57]  = A[1][4][57] ^ D[1][57];
    assign A_theta[1][4][58]  = A[1][4][58] ^ D[1][58];
    assign A_theta[1][4][59]  = A[1][4][59] ^ D[1][59];
    assign A_theta[1][4][60]  = A[1][4][60] ^ D[1][60];
    assign A_theta[1][4][61]  = A[1][4][61] ^ D[1][61];
    assign A_theta[1][4][62]  = A[1][4][62] ^ D[1][62];
    assign A_theta[1][4][63]  = A[1][4][63] ^ D[1][63];
    assign A_theta[2][0][0]  = A[2][0][0] ^ D[2][0];
    assign A_theta[2][0][1]  = A[2][0][1] ^ D[2][1];
    assign A_theta[2][0][2]  = A[2][0][2] ^ D[2][2];
    assign A_theta[2][0][3]  = A[2][0][3] ^ D[2][3];
    assign A_theta[2][0][4]  = A[2][0][4] ^ D[2][4];
    assign A_theta[2][0][5]  = A[2][0][5] ^ D[2][5];
    assign A_theta[2][0][6]  = A[2][0][6] ^ D[2][6];
    assign A_theta[2][0][7]  = A[2][0][7] ^ D[2][7];
    assign A_theta[2][0][8]  = A[2][0][8] ^ D[2][8];
    assign A_theta[2][0][9]  = A[2][0][9] ^ D[2][9];
    assign A_theta[2][0][10]  = A[2][0][10] ^ D[2][10];
    assign A_theta[2][0][11]  = A[2][0][11] ^ D[2][11];
    assign A_theta[2][0][12]  = A[2][0][12] ^ D[2][12];
    assign A_theta[2][0][13]  = A[2][0][13] ^ D[2][13];
    assign A_theta[2][0][14]  = A[2][0][14] ^ D[2][14];
    assign A_theta[2][0][15]  = A[2][0][15] ^ D[2][15];
    assign A_theta[2][0][16]  = A[2][0][16] ^ D[2][16];
    assign A_theta[2][0][17]  = A[2][0][17] ^ D[2][17];
    assign A_theta[2][0][18]  = A[2][0][18] ^ D[2][18];
    assign A_theta[2][0][19]  = A[2][0][19] ^ D[2][19];
    assign A_theta[2][0][20]  = A[2][0][20] ^ D[2][20];
    assign A_theta[2][0][21]  = A[2][0][21] ^ D[2][21];
    assign A_theta[2][0][22]  = A[2][0][22] ^ D[2][22];
    assign A_theta[2][0][23]  = A[2][0][23] ^ D[2][23];
    assign A_theta[2][0][24]  = A[2][0][24] ^ D[2][24];
    assign A_theta[2][0][25]  = A[2][0][25] ^ D[2][25];
    assign A_theta[2][0][26]  = A[2][0][26] ^ D[2][26];
    assign A_theta[2][0][27]  = A[2][0][27] ^ D[2][27];
    assign A_theta[2][0][28]  = A[2][0][28] ^ D[2][28];
    assign A_theta[2][0][29]  = A[2][0][29] ^ D[2][29];
    assign A_theta[2][0][30]  = A[2][0][30] ^ D[2][30];
    assign A_theta[2][0][31]  = A[2][0][31] ^ D[2][31];
    assign A_theta[2][0][32]  = A[2][0][32] ^ D[2][32];
    assign A_theta[2][0][33]  = A[2][0][33] ^ D[2][33];
    assign A_theta[2][0][34]  = A[2][0][34] ^ D[2][34];
    assign A_theta[2][0][35]  = A[2][0][35] ^ D[2][35];
    assign A_theta[2][0][36]  = A[2][0][36] ^ D[2][36];
    assign A_theta[2][0][37]  = A[2][0][37] ^ D[2][37];
    assign A_theta[2][0][38]  = A[2][0][38] ^ D[2][38];
    assign A_theta[2][0][39]  = A[2][0][39] ^ D[2][39];
    assign A_theta[2][0][40]  = A[2][0][40] ^ D[2][40];
    assign A_theta[2][0][41]  = A[2][0][41] ^ D[2][41];
    assign A_theta[2][0][42]  = A[2][0][42] ^ D[2][42];
    assign A_theta[2][0][43]  = A[2][0][43] ^ D[2][43];
    assign A_theta[2][0][44]  = A[2][0][44] ^ D[2][44];
    assign A_theta[2][0][45]  = A[2][0][45] ^ D[2][45];
    assign A_theta[2][0][46]  = A[2][0][46] ^ D[2][46];
    assign A_theta[2][0][47]  = A[2][0][47] ^ D[2][47];
    assign A_theta[2][0][48]  = A[2][0][48] ^ D[2][48];
    assign A_theta[2][0][49]  = A[2][0][49] ^ D[2][49];
    assign A_theta[2][0][50]  = A[2][0][50] ^ D[2][50];
    assign A_theta[2][0][51]  = A[2][0][51] ^ D[2][51];
    assign A_theta[2][0][52]  = A[2][0][52] ^ D[2][52];
    assign A_theta[2][0][53]  = A[2][0][53] ^ D[2][53];
    assign A_theta[2][0][54]  = A[2][0][54] ^ D[2][54];
    assign A_theta[2][0][55]  = A[2][0][55] ^ D[2][55];
    assign A_theta[2][0][56]  = A[2][0][56] ^ D[2][56];
    assign A_theta[2][0][57]  = A[2][0][57] ^ D[2][57];
    assign A_theta[2][0][58]  = A[2][0][58] ^ D[2][58];
    assign A_theta[2][0][59]  = A[2][0][59] ^ D[2][59];
    assign A_theta[2][0][60]  = A[2][0][60] ^ D[2][60];
    assign A_theta[2][0][61]  = A[2][0][61] ^ D[2][61];
    assign A_theta[2][0][62]  = A[2][0][62] ^ D[2][62];
    assign A_theta[2][0][63]  = A[2][0][63] ^ D[2][63];
    assign A_theta[2][1][0]  = A[2][1][0] ^ D[2][0];
    assign A_theta[2][1][1]  = A[2][1][1] ^ D[2][1];
    assign A_theta[2][1][2]  = A[2][1][2] ^ D[2][2];
    assign A_theta[2][1][3]  = A[2][1][3] ^ D[2][3];
    assign A_theta[2][1][4]  = A[2][1][4] ^ D[2][4];
    assign A_theta[2][1][5]  = A[2][1][5] ^ D[2][5];
    assign A_theta[2][1][6]  = A[2][1][6] ^ D[2][6];
    assign A_theta[2][1][7]  = A[2][1][7] ^ D[2][7];
    assign A_theta[2][1][8]  = A[2][1][8] ^ D[2][8];
    assign A_theta[2][1][9]  = A[2][1][9] ^ D[2][9];
    assign A_theta[2][1][10]  = A[2][1][10] ^ D[2][10];
    assign A_theta[2][1][11]  = A[2][1][11] ^ D[2][11];
    assign A_theta[2][1][12]  = A[2][1][12] ^ D[2][12];
    assign A_theta[2][1][13]  = A[2][1][13] ^ D[2][13];
    assign A_theta[2][1][14]  = A[2][1][14] ^ D[2][14];
    assign A_theta[2][1][15]  = A[2][1][15] ^ D[2][15];
    assign A_theta[2][1][16]  = A[2][1][16] ^ D[2][16];
    assign A_theta[2][1][17]  = A[2][1][17] ^ D[2][17];
    assign A_theta[2][1][18]  = A[2][1][18] ^ D[2][18];
    assign A_theta[2][1][19]  = A[2][1][19] ^ D[2][19];
    assign A_theta[2][1][20]  = A[2][1][20] ^ D[2][20];
    assign A_theta[2][1][21]  = A[2][1][21] ^ D[2][21];
    assign A_theta[2][1][22]  = A[2][1][22] ^ D[2][22];
    assign A_theta[2][1][23]  = A[2][1][23] ^ D[2][23];
    assign A_theta[2][1][24]  = A[2][1][24] ^ D[2][24];
    assign A_theta[2][1][25]  = A[2][1][25] ^ D[2][25];
    assign A_theta[2][1][26]  = A[2][1][26] ^ D[2][26];
    assign A_theta[2][1][27]  = A[2][1][27] ^ D[2][27];
    assign A_theta[2][1][28]  = A[2][1][28] ^ D[2][28];
    assign A_theta[2][1][29]  = A[2][1][29] ^ D[2][29];
    assign A_theta[2][1][30]  = A[2][1][30] ^ D[2][30];
    assign A_theta[2][1][31]  = A[2][1][31] ^ D[2][31];
    assign A_theta[2][1][32]  = A[2][1][32] ^ D[2][32];
    assign A_theta[2][1][33]  = A[2][1][33] ^ D[2][33];
    assign A_theta[2][1][34]  = A[2][1][34] ^ D[2][34];
    assign A_theta[2][1][35]  = A[2][1][35] ^ D[2][35];
    assign A_theta[2][1][36]  = A[2][1][36] ^ D[2][36];
    assign A_theta[2][1][37]  = A[2][1][37] ^ D[2][37];
    assign A_theta[2][1][38]  = A[2][1][38] ^ D[2][38];
    assign A_theta[2][1][39]  = A[2][1][39] ^ D[2][39];
    assign A_theta[2][1][40]  = A[2][1][40] ^ D[2][40];
    assign A_theta[2][1][41]  = A[2][1][41] ^ D[2][41];
    assign A_theta[2][1][42]  = A[2][1][42] ^ D[2][42];
    assign A_theta[2][1][43]  = A[2][1][43] ^ D[2][43];
    assign A_theta[2][1][44]  = A[2][1][44] ^ D[2][44];
    assign A_theta[2][1][45]  = A[2][1][45] ^ D[2][45];
    assign A_theta[2][1][46]  = A[2][1][46] ^ D[2][46];
    assign A_theta[2][1][47]  = A[2][1][47] ^ D[2][47];
    assign A_theta[2][1][48]  = A[2][1][48] ^ D[2][48];
    assign A_theta[2][1][49]  = A[2][1][49] ^ D[2][49];
    assign A_theta[2][1][50]  = A[2][1][50] ^ D[2][50];
    assign A_theta[2][1][51]  = A[2][1][51] ^ D[2][51];
    assign A_theta[2][1][52]  = A[2][1][52] ^ D[2][52];
    assign A_theta[2][1][53]  = A[2][1][53] ^ D[2][53];
    assign A_theta[2][1][54]  = A[2][1][54] ^ D[2][54];
    assign A_theta[2][1][55]  = A[2][1][55] ^ D[2][55];
    assign A_theta[2][1][56]  = A[2][1][56] ^ D[2][56];
    assign A_theta[2][1][57]  = A[2][1][57] ^ D[2][57];
    assign A_theta[2][1][58]  = A[2][1][58] ^ D[2][58];
    assign A_theta[2][1][59]  = A[2][1][59] ^ D[2][59];
    assign A_theta[2][1][60]  = A[2][1][60] ^ D[2][60];
    assign A_theta[2][1][61]  = A[2][1][61] ^ D[2][61];
    assign A_theta[2][1][62]  = A[2][1][62] ^ D[2][62];
    assign A_theta[2][1][63]  = A[2][1][63] ^ D[2][63];
    assign A_theta[2][2][0]  = A[2][2][0] ^ D[2][0];
    assign A_theta[2][2][1]  = A[2][2][1] ^ D[2][1];
    assign A_theta[2][2][2]  = A[2][2][2] ^ D[2][2];
    assign A_theta[2][2][3]  = A[2][2][3] ^ D[2][3];
    assign A_theta[2][2][4]  = A[2][2][4] ^ D[2][4];
    assign A_theta[2][2][5]  = A[2][2][5] ^ D[2][5];
    assign A_theta[2][2][6]  = A[2][2][6] ^ D[2][6];
    assign A_theta[2][2][7]  = A[2][2][7] ^ D[2][7];
    assign A_theta[2][2][8]  = A[2][2][8] ^ D[2][8];
    assign A_theta[2][2][9]  = A[2][2][9] ^ D[2][9];
    assign A_theta[2][2][10]  = A[2][2][10] ^ D[2][10];
    assign A_theta[2][2][11]  = A[2][2][11] ^ D[2][11];
    assign A_theta[2][2][12]  = A[2][2][12] ^ D[2][12];
    assign A_theta[2][2][13]  = A[2][2][13] ^ D[2][13];
    assign A_theta[2][2][14]  = A[2][2][14] ^ D[2][14];
    assign A_theta[2][2][15]  = A[2][2][15] ^ D[2][15];
    assign A_theta[2][2][16]  = A[2][2][16] ^ D[2][16];
    assign A_theta[2][2][17]  = A[2][2][17] ^ D[2][17];
    assign A_theta[2][2][18]  = A[2][2][18] ^ D[2][18];
    assign A_theta[2][2][19]  = A[2][2][19] ^ D[2][19];
    assign A_theta[2][2][20]  = A[2][2][20] ^ D[2][20];
    assign A_theta[2][2][21]  = A[2][2][21] ^ D[2][21];
    assign A_theta[2][2][22]  = A[2][2][22] ^ D[2][22];
    assign A_theta[2][2][23]  = A[2][2][23] ^ D[2][23];
    assign A_theta[2][2][24]  = A[2][2][24] ^ D[2][24];
    assign A_theta[2][2][25]  = A[2][2][25] ^ D[2][25];
    assign A_theta[2][2][26]  = A[2][2][26] ^ D[2][26];
    assign A_theta[2][2][27]  = A[2][2][27] ^ D[2][27];
    assign A_theta[2][2][28]  = A[2][2][28] ^ D[2][28];
    assign A_theta[2][2][29]  = A[2][2][29] ^ D[2][29];
    assign A_theta[2][2][30]  = A[2][2][30] ^ D[2][30];
    assign A_theta[2][2][31]  = A[2][2][31] ^ D[2][31];
    assign A_theta[2][2][32]  = A[2][2][32] ^ D[2][32];
    assign A_theta[2][2][33]  = A[2][2][33] ^ D[2][33];
    assign A_theta[2][2][34]  = A[2][2][34] ^ D[2][34];
    assign A_theta[2][2][35]  = A[2][2][35] ^ D[2][35];
    assign A_theta[2][2][36]  = A[2][2][36] ^ D[2][36];
    assign A_theta[2][2][37]  = A[2][2][37] ^ D[2][37];
    assign A_theta[2][2][38]  = A[2][2][38] ^ D[2][38];
    assign A_theta[2][2][39]  = A[2][2][39] ^ D[2][39];
    assign A_theta[2][2][40]  = A[2][2][40] ^ D[2][40];
    assign A_theta[2][2][41]  = A[2][2][41] ^ D[2][41];
    assign A_theta[2][2][42]  = A[2][2][42] ^ D[2][42];
    assign A_theta[2][2][43]  = A[2][2][43] ^ D[2][43];
    assign A_theta[2][2][44]  = A[2][2][44] ^ D[2][44];
    assign A_theta[2][2][45]  = A[2][2][45] ^ D[2][45];
    assign A_theta[2][2][46]  = A[2][2][46] ^ D[2][46];
    assign A_theta[2][2][47]  = A[2][2][47] ^ D[2][47];
    assign A_theta[2][2][48]  = A[2][2][48] ^ D[2][48];
    assign A_theta[2][2][49]  = A[2][2][49] ^ D[2][49];
    assign A_theta[2][2][50]  = A[2][2][50] ^ D[2][50];
    assign A_theta[2][2][51]  = A[2][2][51] ^ D[2][51];
    assign A_theta[2][2][52]  = A[2][2][52] ^ D[2][52];
    assign A_theta[2][2][53]  = A[2][2][53] ^ D[2][53];
    assign A_theta[2][2][54]  = A[2][2][54] ^ D[2][54];
    assign A_theta[2][2][55]  = A[2][2][55] ^ D[2][55];
    assign A_theta[2][2][56]  = A[2][2][56] ^ D[2][56];
    assign A_theta[2][2][57]  = A[2][2][57] ^ D[2][57];
    assign A_theta[2][2][58]  = A[2][2][58] ^ D[2][58];
    assign A_theta[2][2][59]  = A[2][2][59] ^ D[2][59];
    assign A_theta[2][2][60]  = A[2][2][60] ^ D[2][60];
    assign A_theta[2][2][61]  = A[2][2][61] ^ D[2][61];
    assign A_theta[2][2][62]  = A[2][2][62] ^ D[2][62];
    assign A_theta[2][2][63]  = A[2][2][63] ^ D[2][63];
    assign A_theta[2][3][0]  = A[2][3][0] ^ D[2][0];
    assign A_theta[2][3][1]  = A[2][3][1] ^ D[2][1];
    assign A_theta[2][3][2]  = A[2][3][2] ^ D[2][2];
    assign A_theta[2][3][3]  = A[2][3][3] ^ D[2][3];
    assign A_theta[2][3][4]  = A[2][3][4] ^ D[2][4];
    assign A_theta[2][3][5]  = A[2][3][5] ^ D[2][5];
    assign A_theta[2][3][6]  = A[2][3][6] ^ D[2][6];
    assign A_theta[2][3][7]  = A[2][3][7] ^ D[2][7];
    assign A_theta[2][3][8]  = A[2][3][8] ^ D[2][8];
    assign A_theta[2][3][9]  = A[2][3][9] ^ D[2][9];
    assign A_theta[2][3][10]  = A[2][3][10] ^ D[2][10];
    assign A_theta[2][3][11]  = A[2][3][11] ^ D[2][11];
    assign A_theta[2][3][12]  = A[2][3][12] ^ D[2][12];
    assign A_theta[2][3][13]  = A[2][3][13] ^ D[2][13];
    assign A_theta[2][3][14]  = A[2][3][14] ^ D[2][14];
    assign A_theta[2][3][15]  = A[2][3][15] ^ D[2][15];
    assign A_theta[2][3][16]  = A[2][3][16] ^ D[2][16];
    assign A_theta[2][3][17]  = A[2][3][17] ^ D[2][17];
    assign A_theta[2][3][18]  = A[2][3][18] ^ D[2][18];
    assign A_theta[2][3][19]  = A[2][3][19] ^ D[2][19];
    assign A_theta[2][3][20]  = A[2][3][20] ^ D[2][20];
    assign A_theta[2][3][21]  = A[2][3][21] ^ D[2][21];
    assign A_theta[2][3][22]  = A[2][3][22] ^ D[2][22];
    assign A_theta[2][3][23]  = A[2][3][23] ^ D[2][23];
    assign A_theta[2][3][24]  = A[2][3][24] ^ D[2][24];
    assign A_theta[2][3][25]  = A[2][3][25] ^ D[2][25];
    assign A_theta[2][3][26]  = A[2][3][26] ^ D[2][26];
    assign A_theta[2][3][27]  = A[2][3][27] ^ D[2][27];
    assign A_theta[2][3][28]  = A[2][3][28] ^ D[2][28];
    assign A_theta[2][3][29]  = A[2][3][29] ^ D[2][29];
    assign A_theta[2][3][30]  = A[2][3][30] ^ D[2][30];
    assign A_theta[2][3][31]  = A[2][3][31] ^ D[2][31];
    assign A_theta[2][3][32]  = A[2][3][32] ^ D[2][32];
    assign A_theta[2][3][33]  = A[2][3][33] ^ D[2][33];
    assign A_theta[2][3][34]  = A[2][3][34] ^ D[2][34];
    assign A_theta[2][3][35]  = A[2][3][35] ^ D[2][35];
    assign A_theta[2][3][36]  = A[2][3][36] ^ D[2][36];
    assign A_theta[2][3][37]  = A[2][3][37] ^ D[2][37];
    assign A_theta[2][3][38]  = A[2][3][38] ^ D[2][38];
    assign A_theta[2][3][39]  = A[2][3][39] ^ D[2][39];
    assign A_theta[2][3][40]  = A[2][3][40] ^ D[2][40];
    assign A_theta[2][3][41]  = A[2][3][41] ^ D[2][41];
    assign A_theta[2][3][42]  = A[2][3][42] ^ D[2][42];
    assign A_theta[2][3][43]  = A[2][3][43] ^ D[2][43];
    assign A_theta[2][3][44]  = A[2][3][44] ^ D[2][44];
    assign A_theta[2][3][45]  = A[2][3][45] ^ D[2][45];
    assign A_theta[2][3][46]  = A[2][3][46] ^ D[2][46];
    assign A_theta[2][3][47]  = A[2][3][47] ^ D[2][47];
    assign A_theta[2][3][48]  = A[2][3][48] ^ D[2][48];
    assign A_theta[2][3][49]  = A[2][3][49] ^ D[2][49];
    assign A_theta[2][3][50]  = A[2][3][50] ^ D[2][50];
    assign A_theta[2][3][51]  = A[2][3][51] ^ D[2][51];
    assign A_theta[2][3][52]  = A[2][3][52] ^ D[2][52];
    assign A_theta[2][3][53]  = A[2][3][53] ^ D[2][53];
    assign A_theta[2][3][54]  = A[2][3][54] ^ D[2][54];
    assign A_theta[2][3][55]  = A[2][3][55] ^ D[2][55];
    assign A_theta[2][3][56]  = A[2][3][56] ^ D[2][56];
    assign A_theta[2][3][57]  = A[2][3][57] ^ D[2][57];
    assign A_theta[2][3][58]  = A[2][3][58] ^ D[2][58];
    assign A_theta[2][3][59]  = A[2][3][59] ^ D[2][59];
    assign A_theta[2][3][60]  = A[2][3][60] ^ D[2][60];
    assign A_theta[2][3][61]  = A[2][3][61] ^ D[2][61];
    assign A_theta[2][3][62]  = A[2][3][62] ^ D[2][62];
    assign A_theta[2][3][63]  = A[2][3][63] ^ D[2][63];
    assign A_theta[2][4][0]  = A[2][4][0] ^ D[2][0];
    assign A_theta[2][4][1]  = A[2][4][1] ^ D[2][1];
    assign A_theta[2][4][2]  = A[2][4][2] ^ D[2][2];
    assign A_theta[2][4][3]  = A[2][4][3] ^ D[2][3];
    assign A_theta[2][4][4]  = A[2][4][4] ^ D[2][4];
    assign A_theta[2][4][5]  = A[2][4][5] ^ D[2][5];
    assign A_theta[2][4][6]  = A[2][4][6] ^ D[2][6];
    assign A_theta[2][4][7]  = A[2][4][7] ^ D[2][7];
    assign A_theta[2][4][8]  = A[2][4][8] ^ D[2][8];
    assign A_theta[2][4][9]  = A[2][4][9] ^ D[2][9];
    assign A_theta[2][4][10]  = A[2][4][10] ^ D[2][10];
    assign A_theta[2][4][11]  = A[2][4][11] ^ D[2][11];
    assign A_theta[2][4][12]  = A[2][4][12] ^ D[2][12];
    assign A_theta[2][4][13]  = A[2][4][13] ^ D[2][13];
    assign A_theta[2][4][14]  = A[2][4][14] ^ D[2][14];
    assign A_theta[2][4][15]  = A[2][4][15] ^ D[2][15];
    assign A_theta[2][4][16]  = A[2][4][16] ^ D[2][16];
    assign A_theta[2][4][17]  = A[2][4][17] ^ D[2][17];
    assign A_theta[2][4][18]  = A[2][4][18] ^ D[2][18];
    assign A_theta[2][4][19]  = A[2][4][19] ^ D[2][19];
    assign A_theta[2][4][20]  = A[2][4][20] ^ D[2][20];
    assign A_theta[2][4][21]  = A[2][4][21] ^ D[2][21];
    assign A_theta[2][4][22]  = A[2][4][22] ^ D[2][22];
    assign A_theta[2][4][23]  = A[2][4][23] ^ D[2][23];
    assign A_theta[2][4][24]  = A[2][4][24] ^ D[2][24];
    assign A_theta[2][4][25]  = A[2][4][25] ^ D[2][25];
    assign A_theta[2][4][26]  = A[2][4][26] ^ D[2][26];
    assign A_theta[2][4][27]  = A[2][4][27] ^ D[2][27];
    assign A_theta[2][4][28]  = A[2][4][28] ^ D[2][28];
    assign A_theta[2][4][29]  = A[2][4][29] ^ D[2][29];
    assign A_theta[2][4][30]  = A[2][4][30] ^ D[2][30];
    assign A_theta[2][4][31]  = A[2][4][31] ^ D[2][31];
    assign A_theta[2][4][32]  = A[2][4][32] ^ D[2][32];
    assign A_theta[2][4][33]  = A[2][4][33] ^ D[2][33];
    assign A_theta[2][4][34]  = A[2][4][34] ^ D[2][34];
    assign A_theta[2][4][35]  = A[2][4][35] ^ D[2][35];
    assign A_theta[2][4][36]  = A[2][4][36] ^ D[2][36];
    assign A_theta[2][4][37]  = A[2][4][37] ^ D[2][37];
    assign A_theta[2][4][38]  = A[2][4][38] ^ D[2][38];
    assign A_theta[2][4][39]  = A[2][4][39] ^ D[2][39];
    assign A_theta[2][4][40]  = A[2][4][40] ^ D[2][40];
    assign A_theta[2][4][41]  = A[2][4][41] ^ D[2][41];
    assign A_theta[2][4][42]  = A[2][4][42] ^ D[2][42];
    assign A_theta[2][4][43]  = A[2][4][43] ^ D[2][43];
    assign A_theta[2][4][44]  = A[2][4][44] ^ D[2][44];
    assign A_theta[2][4][45]  = A[2][4][45] ^ D[2][45];
    assign A_theta[2][4][46]  = A[2][4][46] ^ D[2][46];
    assign A_theta[2][4][47]  = A[2][4][47] ^ D[2][47];
    assign A_theta[2][4][48]  = A[2][4][48] ^ D[2][48];
    assign A_theta[2][4][49]  = A[2][4][49] ^ D[2][49];
    assign A_theta[2][4][50]  = A[2][4][50] ^ D[2][50];
    assign A_theta[2][4][51]  = A[2][4][51] ^ D[2][51];
    assign A_theta[2][4][52]  = A[2][4][52] ^ D[2][52];
    assign A_theta[2][4][53]  = A[2][4][53] ^ D[2][53];
    assign A_theta[2][4][54]  = A[2][4][54] ^ D[2][54];
    assign A_theta[2][4][55]  = A[2][4][55] ^ D[2][55];
    assign A_theta[2][4][56]  = A[2][4][56] ^ D[2][56];
    assign A_theta[2][4][57]  = A[2][4][57] ^ D[2][57];
    assign A_theta[2][4][58]  = A[2][4][58] ^ D[2][58];
    assign A_theta[2][4][59]  = A[2][4][59] ^ D[2][59];
    assign A_theta[2][4][60]  = A[2][4][60] ^ D[2][60];
    assign A_theta[2][4][61]  = A[2][4][61] ^ D[2][61];
    assign A_theta[2][4][62]  = A[2][4][62] ^ D[2][62];
    assign A_theta[2][4][63]  = A[2][4][63] ^ D[2][63];
    assign A_theta[3][0][0]  = A[3][0][0] ^ D[3][0];
    assign A_theta[3][0][1]  = A[3][0][1] ^ D[3][1];
    assign A_theta[3][0][2]  = A[3][0][2] ^ D[3][2];
    assign A_theta[3][0][3]  = A[3][0][3] ^ D[3][3];
    assign A_theta[3][0][4]  = A[3][0][4] ^ D[3][4];
    assign A_theta[3][0][5]  = A[3][0][5] ^ D[3][5];
    assign A_theta[3][0][6]  = A[3][0][6] ^ D[3][6];
    assign A_theta[3][0][7]  = A[3][0][7] ^ D[3][7];
    assign A_theta[3][0][8]  = A[3][0][8] ^ D[3][8];
    assign A_theta[3][0][9]  = A[3][0][9] ^ D[3][9];
    assign A_theta[3][0][10]  = A[3][0][10] ^ D[3][10];
    assign A_theta[3][0][11]  = A[3][0][11] ^ D[3][11];
    assign A_theta[3][0][12]  = A[3][0][12] ^ D[3][12];
    assign A_theta[3][0][13]  = A[3][0][13] ^ D[3][13];
    assign A_theta[3][0][14]  = A[3][0][14] ^ D[3][14];
    assign A_theta[3][0][15]  = A[3][0][15] ^ D[3][15];
    assign A_theta[3][0][16]  = A[3][0][16] ^ D[3][16];
    assign A_theta[3][0][17]  = A[3][0][17] ^ D[3][17];
    assign A_theta[3][0][18]  = A[3][0][18] ^ D[3][18];
    assign A_theta[3][0][19]  = A[3][0][19] ^ D[3][19];
    assign A_theta[3][0][20]  = A[3][0][20] ^ D[3][20];
    assign A_theta[3][0][21]  = A[3][0][21] ^ D[3][21];
    assign A_theta[3][0][22]  = A[3][0][22] ^ D[3][22];
    assign A_theta[3][0][23]  = A[3][0][23] ^ D[3][23];
    assign A_theta[3][0][24]  = A[3][0][24] ^ D[3][24];
    assign A_theta[3][0][25]  = A[3][0][25] ^ D[3][25];
    assign A_theta[3][0][26]  = A[3][0][26] ^ D[3][26];
    assign A_theta[3][0][27]  = A[3][0][27] ^ D[3][27];
    assign A_theta[3][0][28]  = A[3][0][28] ^ D[3][28];
    assign A_theta[3][0][29]  = A[3][0][29] ^ D[3][29];
    assign A_theta[3][0][30]  = A[3][0][30] ^ D[3][30];
    assign A_theta[3][0][31]  = A[3][0][31] ^ D[3][31];
    assign A_theta[3][0][32]  = A[3][0][32] ^ D[3][32];
    assign A_theta[3][0][33]  = A[3][0][33] ^ D[3][33];
    assign A_theta[3][0][34]  = A[3][0][34] ^ D[3][34];
    assign A_theta[3][0][35]  = A[3][0][35] ^ D[3][35];
    assign A_theta[3][0][36]  = A[3][0][36] ^ D[3][36];
    assign A_theta[3][0][37]  = A[3][0][37] ^ D[3][37];
    assign A_theta[3][0][38]  = A[3][0][38] ^ D[3][38];
    assign A_theta[3][0][39]  = A[3][0][39] ^ D[3][39];
    assign A_theta[3][0][40]  = A[3][0][40] ^ D[3][40];
    assign A_theta[3][0][41]  = A[3][0][41] ^ D[3][41];
    assign A_theta[3][0][42]  = A[3][0][42] ^ D[3][42];
    assign A_theta[3][0][43]  = A[3][0][43] ^ D[3][43];
    assign A_theta[3][0][44]  = A[3][0][44] ^ D[3][44];
    assign A_theta[3][0][45]  = A[3][0][45] ^ D[3][45];
    assign A_theta[3][0][46]  = A[3][0][46] ^ D[3][46];
    assign A_theta[3][0][47]  = A[3][0][47] ^ D[3][47];
    assign A_theta[3][0][48]  = A[3][0][48] ^ D[3][48];
    assign A_theta[3][0][49]  = A[3][0][49] ^ D[3][49];
    assign A_theta[3][0][50]  = A[3][0][50] ^ D[3][50];
    assign A_theta[3][0][51]  = A[3][0][51] ^ D[3][51];
    assign A_theta[3][0][52]  = A[3][0][52] ^ D[3][52];
    assign A_theta[3][0][53]  = A[3][0][53] ^ D[3][53];
    assign A_theta[3][0][54]  = A[3][0][54] ^ D[3][54];
    assign A_theta[3][0][55]  = A[3][0][55] ^ D[3][55];
    assign A_theta[3][0][56]  = A[3][0][56] ^ D[3][56];
    assign A_theta[3][0][57]  = A[3][0][57] ^ D[3][57];
    assign A_theta[3][0][58]  = A[3][0][58] ^ D[3][58];
    assign A_theta[3][0][59]  = A[3][0][59] ^ D[3][59];
    assign A_theta[3][0][60]  = A[3][0][60] ^ D[3][60];
    assign A_theta[3][0][61]  = A[3][0][61] ^ D[3][61];
    assign A_theta[3][0][62]  = A[3][0][62] ^ D[3][62];
    assign A_theta[3][0][63]  = A[3][0][63] ^ D[3][63];
    assign A_theta[3][1][0]  = A[3][1][0] ^ D[3][0];
    assign A_theta[3][1][1]  = A[3][1][1] ^ D[3][1];
    assign A_theta[3][1][2]  = A[3][1][2] ^ D[3][2];
    assign A_theta[3][1][3]  = A[3][1][3] ^ D[3][3];
    assign A_theta[3][1][4]  = A[3][1][4] ^ D[3][4];
    assign A_theta[3][1][5]  = A[3][1][5] ^ D[3][5];
    assign A_theta[3][1][6]  = A[3][1][6] ^ D[3][6];
    assign A_theta[3][1][7]  = A[3][1][7] ^ D[3][7];
    assign A_theta[3][1][8]  = A[3][1][8] ^ D[3][8];
    assign A_theta[3][1][9]  = A[3][1][9] ^ D[3][9];
    assign A_theta[3][1][10]  = A[3][1][10] ^ D[3][10];
    assign A_theta[3][1][11]  = A[3][1][11] ^ D[3][11];
    assign A_theta[3][1][12]  = A[3][1][12] ^ D[3][12];
    assign A_theta[3][1][13]  = A[3][1][13] ^ D[3][13];
    assign A_theta[3][1][14]  = A[3][1][14] ^ D[3][14];
    assign A_theta[3][1][15]  = A[3][1][15] ^ D[3][15];
    assign A_theta[3][1][16]  = A[3][1][16] ^ D[3][16];
    assign A_theta[3][1][17]  = A[3][1][17] ^ D[3][17];
    assign A_theta[3][1][18]  = A[3][1][18] ^ D[3][18];
    assign A_theta[3][1][19]  = A[3][1][19] ^ D[3][19];
    assign A_theta[3][1][20]  = A[3][1][20] ^ D[3][20];
    assign A_theta[3][1][21]  = A[3][1][21] ^ D[3][21];
    assign A_theta[3][1][22]  = A[3][1][22] ^ D[3][22];
    assign A_theta[3][1][23]  = A[3][1][23] ^ D[3][23];
    assign A_theta[3][1][24]  = A[3][1][24] ^ D[3][24];
    assign A_theta[3][1][25]  = A[3][1][25] ^ D[3][25];
    assign A_theta[3][1][26]  = A[3][1][26] ^ D[3][26];
    assign A_theta[3][1][27]  = A[3][1][27] ^ D[3][27];
    assign A_theta[3][1][28]  = A[3][1][28] ^ D[3][28];
    assign A_theta[3][1][29]  = A[3][1][29] ^ D[3][29];
    assign A_theta[3][1][30]  = A[3][1][30] ^ D[3][30];
    assign A_theta[3][1][31]  = A[3][1][31] ^ D[3][31];
    assign A_theta[3][1][32]  = A[3][1][32] ^ D[3][32];
    assign A_theta[3][1][33]  = A[3][1][33] ^ D[3][33];
    assign A_theta[3][1][34]  = A[3][1][34] ^ D[3][34];
    assign A_theta[3][1][35]  = A[3][1][35] ^ D[3][35];
    assign A_theta[3][1][36]  = A[3][1][36] ^ D[3][36];
    assign A_theta[3][1][37]  = A[3][1][37] ^ D[3][37];
    assign A_theta[3][1][38]  = A[3][1][38] ^ D[3][38];
    assign A_theta[3][1][39]  = A[3][1][39] ^ D[3][39];
    assign A_theta[3][1][40]  = A[3][1][40] ^ D[3][40];
    assign A_theta[3][1][41]  = A[3][1][41] ^ D[3][41];
    assign A_theta[3][1][42]  = A[3][1][42] ^ D[3][42];
    assign A_theta[3][1][43]  = A[3][1][43] ^ D[3][43];
    assign A_theta[3][1][44]  = A[3][1][44] ^ D[3][44];
    assign A_theta[3][1][45]  = A[3][1][45] ^ D[3][45];
    assign A_theta[3][1][46]  = A[3][1][46] ^ D[3][46];
    assign A_theta[3][1][47]  = A[3][1][47] ^ D[3][47];
    assign A_theta[3][1][48]  = A[3][1][48] ^ D[3][48];
    assign A_theta[3][1][49]  = A[3][1][49] ^ D[3][49];
    assign A_theta[3][1][50]  = A[3][1][50] ^ D[3][50];
    assign A_theta[3][1][51]  = A[3][1][51] ^ D[3][51];
    assign A_theta[3][1][52]  = A[3][1][52] ^ D[3][52];
    assign A_theta[3][1][53]  = A[3][1][53] ^ D[3][53];
    assign A_theta[3][1][54]  = A[3][1][54] ^ D[3][54];
    assign A_theta[3][1][55]  = A[3][1][55] ^ D[3][55];
    assign A_theta[3][1][56]  = A[3][1][56] ^ D[3][56];
    assign A_theta[3][1][57]  = A[3][1][57] ^ D[3][57];
    assign A_theta[3][1][58]  = A[3][1][58] ^ D[3][58];
    assign A_theta[3][1][59]  = A[3][1][59] ^ D[3][59];
    assign A_theta[3][1][60]  = A[3][1][60] ^ D[3][60];
    assign A_theta[3][1][61]  = A[3][1][61] ^ D[3][61];
    assign A_theta[3][1][62]  = A[3][1][62] ^ D[3][62];
    assign A_theta[3][1][63]  = A[3][1][63] ^ D[3][63];
    assign A_theta[3][2][0]  = A[3][2][0] ^ D[3][0];
    assign A_theta[3][2][1]  = A[3][2][1] ^ D[3][1];
    assign A_theta[3][2][2]  = A[3][2][2] ^ D[3][2];
    assign A_theta[3][2][3]  = A[3][2][3] ^ D[3][3];
    assign A_theta[3][2][4]  = A[3][2][4] ^ D[3][4];
    assign A_theta[3][2][5]  = A[3][2][5] ^ D[3][5];
    assign A_theta[3][2][6]  = A[3][2][6] ^ D[3][6];
    assign A_theta[3][2][7]  = A[3][2][7] ^ D[3][7];
    assign A_theta[3][2][8]  = A[3][2][8] ^ D[3][8];
    assign A_theta[3][2][9]  = A[3][2][9] ^ D[3][9];
    assign A_theta[3][2][10]  = A[3][2][10] ^ D[3][10];
    assign A_theta[3][2][11]  = A[3][2][11] ^ D[3][11];
    assign A_theta[3][2][12]  = A[3][2][12] ^ D[3][12];
    assign A_theta[3][2][13]  = A[3][2][13] ^ D[3][13];
    assign A_theta[3][2][14]  = A[3][2][14] ^ D[3][14];
    assign A_theta[3][2][15]  = A[3][2][15] ^ D[3][15];
    assign A_theta[3][2][16]  = A[3][2][16] ^ D[3][16];
    assign A_theta[3][2][17]  = A[3][2][17] ^ D[3][17];
    assign A_theta[3][2][18]  = A[3][2][18] ^ D[3][18];
    assign A_theta[3][2][19]  = A[3][2][19] ^ D[3][19];
    assign A_theta[3][2][20]  = A[3][2][20] ^ D[3][20];
    assign A_theta[3][2][21]  = A[3][2][21] ^ D[3][21];
    assign A_theta[3][2][22]  = A[3][2][22] ^ D[3][22];
    assign A_theta[3][2][23]  = A[3][2][23] ^ D[3][23];
    assign A_theta[3][2][24]  = A[3][2][24] ^ D[3][24];
    assign A_theta[3][2][25]  = A[3][2][25] ^ D[3][25];
    assign A_theta[3][2][26]  = A[3][2][26] ^ D[3][26];
    assign A_theta[3][2][27]  = A[3][2][27] ^ D[3][27];
    assign A_theta[3][2][28]  = A[3][2][28] ^ D[3][28];
    assign A_theta[3][2][29]  = A[3][2][29] ^ D[3][29];
    assign A_theta[3][2][30]  = A[3][2][30] ^ D[3][30];
    assign A_theta[3][2][31]  = A[3][2][31] ^ D[3][31];
    assign A_theta[3][2][32]  = A[3][2][32] ^ D[3][32];
    assign A_theta[3][2][33]  = A[3][2][33] ^ D[3][33];
    assign A_theta[3][2][34]  = A[3][2][34] ^ D[3][34];
    assign A_theta[3][2][35]  = A[3][2][35] ^ D[3][35];
    assign A_theta[3][2][36]  = A[3][2][36] ^ D[3][36];
    assign A_theta[3][2][37]  = A[3][2][37] ^ D[3][37];
    assign A_theta[3][2][38]  = A[3][2][38] ^ D[3][38];
    assign A_theta[3][2][39]  = A[3][2][39] ^ D[3][39];
    assign A_theta[3][2][40]  = A[3][2][40] ^ D[3][40];
    assign A_theta[3][2][41]  = A[3][2][41] ^ D[3][41];
    assign A_theta[3][2][42]  = A[3][2][42] ^ D[3][42];
    assign A_theta[3][2][43]  = A[3][2][43] ^ D[3][43];
    assign A_theta[3][2][44]  = A[3][2][44] ^ D[3][44];
    assign A_theta[3][2][45]  = A[3][2][45] ^ D[3][45];
    assign A_theta[3][2][46]  = A[3][2][46] ^ D[3][46];
    assign A_theta[3][2][47]  = A[3][2][47] ^ D[3][47];
    assign A_theta[3][2][48]  = A[3][2][48] ^ D[3][48];
    assign A_theta[3][2][49]  = A[3][2][49] ^ D[3][49];
    assign A_theta[3][2][50]  = A[3][2][50] ^ D[3][50];
    assign A_theta[3][2][51]  = A[3][2][51] ^ D[3][51];
    assign A_theta[3][2][52]  = A[3][2][52] ^ D[3][52];
    assign A_theta[3][2][53]  = A[3][2][53] ^ D[3][53];
    assign A_theta[3][2][54]  = A[3][2][54] ^ D[3][54];
    assign A_theta[3][2][55]  = A[3][2][55] ^ D[3][55];
    assign A_theta[3][2][56]  = A[3][2][56] ^ D[3][56];
    assign A_theta[3][2][57]  = A[3][2][57] ^ D[3][57];
    assign A_theta[3][2][58]  = A[3][2][58] ^ D[3][58];
    assign A_theta[3][2][59]  = A[3][2][59] ^ D[3][59];
    assign A_theta[3][2][60]  = A[3][2][60] ^ D[3][60];
    assign A_theta[3][2][61]  = A[3][2][61] ^ D[3][61];
    assign A_theta[3][2][62]  = A[3][2][62] ^ D[3][62];
    assign A_theta[3][2][63]  = A[3][2][63] ^ D[3][63];
    assign A_theta[3][3][0]  = A[3][3][0] ^ D[3][0];
    assign A_theta[3][3][1]  = A[3][3][1] ^ D[3][1];
    assign A_theta[3][3][2]  = A[3][3][2] ^ D[3][2];
    assign A_theta[3][3][3]  = A[3][3][3] ^ D[3][3];
    assign A_theta[3][3][4]  = A[3][3][4] ^ D[3][4];
    assign A_theta[3][3][5]  = A[3][3][5] ^ D[3][5];
    assign A_theta[3][3][6]  = A[3][3][6] ^ D[3][6];
    assign A_theta[3][3][7]  = A[3][3][7] ^ D[3][7];
    assign A_theta[3][3][8]  = A[3][3][8] ^ D[3][8];
    assign A_theta[3][3][9]  = A[3][3][9] ^ D[3][9];
    assign A_theta[3][3][10]  = A[3][3][10] ^ D[3][10];
    assign A_theta[3][3][11]  = A[3][3][11] ^ D[3][11];
    assign A_theta[3][3][12]  = A[3][3][12] ^ D[3][12];
    assign A_theta[3][3][13]  = A[3][3][13] ^ D[3][13];
    assign A_theta[3][3][14]  = A[3][3][14] ^ D[3][14];
    assign A_theta[3][3][15]  = A[3][3][15] ^ D[3][15];
    assign A_theta[3][3][16]  = A[3][3][16] ^ D[3][16];
    assign A_theta[3][3][17]  = A[3][3][17] ^ D[3][17];
    assign A_theta[3][3][18]  = A[3][3][18] ^ D[3][18];
    assign A_theta[3][3][19]  = A[3][3][19] ^ D[3][19];
    assign A_theta[3][3][20]  = A[3][3][20] ^ D[3][20];
    assign A_theta[3][3][21]  = A[3][3][21] ^ D[3][21];
    assign A_theta[3][3][22]  = A[3][3][22] ^ D[3][22];
    assign A_theta[3][3][23]  = A[3][3][23] ^ D[3][23];
    assign A_theta[3][3][24]  = A[3][3][24] ^ D[3][24];
    assign A_theta[3][3][25]  = A[3][3][25] ^ D[3][25];
    assign A_theta[3][3][26]  = A[3][3][26] ^ D[3][26];
    assign A_theta[3][3][27]  = A[3][3][27] ^ D[3][27];
    assign A_theta[3][3][28]  = A[3][3][28] ^ D[3][28];
    assign A_theta[3][3][29]  = A[3][3][29] ^ D[3][29];
    assign A_theta[3][3][30]  = A[3][3][30] ^ D[3][30];
    assign A_theta[3][3][31]  = A[3][3][31] ^ D[3][31];
    assign A_theta[3][3][32]  = A[3][3][32] ^ D[3][32];
    assign A_theta[3][3][33]  = A[3][3][33] ^ D[3][33];
    assign A_theta[3][3][34]  = A[3][3][34] ^ D[3][34];
    assign A_theta[3][3][35]  = A[3][3][35] ^ D[3][35];
    assign A_theta[3][3][36]  = A[3][3][36] ^ D[3][36];
    assign A_theta[3][3][37]  = A[3][3][37] ^ D[3][37];
    assign A_theta[3][3][38]  = A[3][3][38] ^ D[3][38];
    assign A_theta[3][3][39]  = A[3][3][39] ^ D[3][39];
    assign A_theta[3][3][40]  = A[3][3][40] ^ D[3][40];
    assign A_theta[3][3][41]  = A[3][3][41] ^ D[3][41];
    assign A_theta[3][3][42]  = A[3][3][42] ^ D[3][42];
    assign A_theta[3][3][43]  = A[3][3][43] ^ D[3][43];
    assign A_theta[3][3][44]  = A[3][3][44] ^ D[3][44];
    assign A_theta[3][3][45]  = A[3][3][45] ^ D[3][45];
    assign A_theta[3][3][46]  = A[3][3][46] ^ D[3][46];
    assign A_theta[3][3][47]  = A[3][3][47] ^ D[3][47];
    assign A_theta[3][3][48]  = A[3][3][48] ^ D[3][48];
    assign A_theta[3][3][49]  = A[3][3][49] ^ D[3][49];
    assign A_theta[3][3][50]  = A[3][3][50] ^ D[3][50];
    assign A_theta[3][3][51]  = A[3][3][51] ^ D[3][51];
    assign A_theta[3][3][52]  = A[3][3][52] ^ D[3][52];
    assign A_theta[3][3][53]  = A[3][3][53] ^ D[3][53];
    assign A_theta[3][3][54]  = A[3][3][54] ^ D[3][54];
    assign A_theta[3][3][55]  = A[3][3][55] ^ D[3][55];
    assign A_theta[3][3][56]  = A[3][3][56] ^ D[3][56];
    assign A_theta[3][3][57]  = A[3][3][57] ^ D[3][57];
    assign A_theta[3][3][58]  = A[3][3][58] ^ D[3][58];
    assign A_theta[3][3][59]  = A[3][3][59] ^ D[3][59];
    assign A_theta[3][3][60]  = A[3][3][60] ^ D[3][60];
    assign A_theta[3][3][61]  = A[3][3][61] ^ D[3][61];
    assign A_theta[3][3][62]  = A[3][3][62] ^ D[3][62];
    assign A_theta[3][3][63]  = A[3][3][63] ^ D[3][63];
    assign A_theta[3][4][0]  = A[3][4][0] ^ D[3][0];
    assign A_theta[3][4][1]  = A[3][4][1] ^ D[3][1];
    assign A_theta[3][4][2]  = A[3][4][2] ^ D[3][2];
    assign A_theta[3][4][3]  = A[3][4][3] ^ D[3][3];
    assign A_theta[3][4][4]  = A[3][4][4] ^ D[3][4];
    assign A_theta[3][4][5]  = A[3][4][5] ^ D[3][5];
    assign A_theta[3][4][6]  = A[3][4][6] ^ D[3][6];
    assign A_theta[3][4][7]  = A[3][4][7] ^ D[3][7];
    assign A_theta[3][4][8]  = A[3][4][8] ^ D[3][8];
    assign A_theta[3][4][9]  = A[3][4][9] ^ D[3][9];
    assign A_theta[3][4][10]  = A[3][4][10] ^ D[3][10];
    assign A_theta[3][4][11]  = A[3][4][11] ^ D[3][11];
    assign A_theta[3][4][12]  = A[3][4][12] ^ D[3][12];
    assign A_theta[3][4][13]  = A[3][4][13] ^ D[3][13];
    assign A_theta[3][4][14]  = A[3][4][14] ^ D[3][14];
    assign A_theta[3][4][15]  = A[3][4][15] ^ D[3][15];
    assign A_theta[3][4][16]  = A[3][4][16] ^ D[3][16];
    assign A_theta[3][4][17]  = A[3][4][17] ^ D[3][17];
    assign A_theta[3][4][18]  = A[3][4][18] ^ D[3][18];
    assign A_theta[3][4][19]  = A[3][4][19] ^ D[3][19];
    assign A_theta[3][4][20]  = A[3][4][20] ^ D[3][20];
    assign A_theta[3][4][21]  = A[3][4][21] ^ D[3][21];
    assign A_theta[3][4][22]  = A[3][4][22] ^ D[3][22];
    assign A_theta[3][4][23]  = A[3][4][23] ^ D[3][23];
    assign A_theta[3][4][24]  = A[3][4][24] ^ D[3][24];
    assign A_theta[3][4][25]  = A[3][4][25] ^ D[3][25];
    assign A_theta[3][4][26]  = A[3][4][26] ^ D[3][26];
    assign A_theta[3][4][27]  = A[3][4][27] ^ D[3][27];
    assign A_theta[3][4][28]  = A[3][4][28] ^ D[3][28];
    assign A_theta[3][4][29]  = A[3][4][29] ^ D[3][29];
    assign A_theta[3][4][30]  = A[3][4][30] ^ D[3][30];
    assign A_theta[3][4][31]  = A[3][4][31] ^ D[3][31];
    assign A_theta[3][4][32]  = A[3][4][32] ^ D[3][32];
    assign A_theta[3][4][33]  = A[3][4][33] ^ D[3][33];
    assign A_theta[3][4][34]  = A[3][4][34] ^ D[3][34];
    assign A_theta[3][4][35]  = A[3][4][35] ^ D[3][35];
    assign A_theta[3][4][36]  = A[3][4][36] ^ D[3][36];
    assign A_theta[3][4][37]  = A[3][4][37] ^ D[3][37];
    assign A_theta[3][4][38]  = A[3][4][38] ^ D[3][38];
    assign A_theta[3][4][39]  = A[3][4][39] ^ D[3][39];
    assign A_theta[3][4][40]  = A[3][4][40] ^ D[3][40];
    assign A_theta[3][4][41]  = A[3][4][41] ^ D[3][41];
    assign A_theta[3][4][42]  = A[3][4][42] ^ D[3][42];
    assign A_theta[3][4][43]  = A[3][4][43] ^ D[3][43];
    assign A_theta[3][4][44]  = A[3][4][44] ^ D[3][44];
    assign A_theta[3][4][45]  = A[3][4][45] ^ D[3][45];
    assign A_theta[3][4][46]  = A[3][4][46] ^ D[3][46];
    assign A_theta[3][4][47]  = A[3][4][47] ^ D[3][47];
    assign A_theta[3][4][48]  = A[3][4][48] ^ D[3][48];
    assign A_theta[3][4][49]  = A[3][4][49] ^ D[3][49];
    assign A_theta[3][4][50]  = A[3][4][50] ^ D[3][50];
    assign A_theta[3][4][51]  = A[3][4][51] ^ D[3][51];
    assign A_theta[3][4][52]  = A[3][4][52] ^ D[3][52];
    assign A_theta[3][4][53]  = A[3][4][53] ^ D[3][53];
    assign A_theta[3][4][54]  = A[3][4][54] ^ D[3][54];
    assign A_theta[3][4][55]  = A[3][4][55] ^ D[3][55];
    assign A_theta[3][4][56]  = A[3][4][56] ^ D[3][56];
    assign A_theta[3][4][57]  = A[3][4][57] ^ D[3][57];
    assign A_theta[3][4][58]  = A[3][4][58] ^ D[3][58];
    assign A_theta[3][4][59]  = A[3][4][59] ^ D[3][59];
    assign A_theta[3][4][60]  = A[3][4][60] ^ D[3][60];
    assign A_theta[3][4][61]  = A[3][4][61] ^ D[3][61];
    assign A_theta[3][4][62]  = A[3][4][62] ^ D[3][62];
    assign A_theta[3][4][63]  = A[3][4][63] ^ D[3][63];
    assign A_theta[4][0][0]  = A[4][0][0] ^ D[4][0];
    assign A_theta[4][0][1]  = A[4][0][1] ^ D[4][1];
    assign A_theta[4][0][2]  = A[4][0][2] ^ D[4][2];
    assign A_theta[4][0][3]  = A[4][0][3] ^ D[4][3];
    assign A_theta[4][0][4]  = A[4][0][4] ^ D[4][4];
    assign A_theta[4][0][5]  = A[4][0][5] ^ D[4][5];
    assign A_theta[4][0][6]  = A[4][0][6] ^ D[4][6];
    assign A_theta[4][0][7]  = A[4][0][7] ^ D[4][7];
    assign A_theta[4][0][8]  = A[4][0][8] ^ D[4][8];
    assign A_theta[4][0][9]  = A[4][0][9] ^ D[4][9];
    assign A_theta[4][0][10]  = A[4][0][10] ^ D[4][10];
    assign A_theta[4][0][11]  = A[4][0][11] ^ D[4][11];
    assign A_theta[4][0][12]  = A[4][0][12] ^ D[4][12];
    assign A_theta[4][0][13]  = A[4][0][13] ^ D[4][13];
    assign A_theta[4][0][14]  = A[4][0][14] ^ D[4][14];
    assign A_theta[4][0][15]  = A[4][0][15] ^ D[4][15];
    assign A_theta[4][0][16]  = A[4][0][16] ^ D[4][16];
    assign A_theta[4][0][17]  = A[4][0][17] ^ D[4][17];
    assign A_theta[4][0][18]  = A[4][0][18] ^ D[4][18];
    assign A_theta[4][0][19]  = A[4][0][19] ^ D[4][19];
    assign A_theta[4][0][20]  = A[4][0][20] ^ D[4][20];
    assign A_theta[4][0][21]  = A[4][0][21] ^ D[4][21];
    assign A_theta[4][0][22]  = A[4][0][22] ^ D[4][22];
    assign A_theta[4][0][23]  = A[4][0][23] ^ D[4][23];
    assign A_theta[4][0][24]  = A[4][0][24] ^ D[4][24];
    assign A_theta[4][0][25]  = A[4][0][25] ^ D[4][25];
    assign A_theta[4][0][26]  = A[4][0][26] ^ D[4][26];
    assign A_theta[4][0][27]  = A[4][0][27] ^ D[4][27];
    assign A_theta[4][0][28]  = A[4][0][28] ^ D[4][28];
    assign A_theta[4][0][29]  = A[4][0][29] ^ D[4][29];
    assign A_theta[4][0][30]  = A[4][0][30] ^ D[4][30];
    assign A_theta[4][0][31]  = A[4][0][31] ^ D[4][31];
    assign A_theta[4][0][32]  = A[4][0][32] ^ D[4][32];
    assign A_theta[4][0][33]  = A[4][0][33] ^ D[4][33];
    assign A_theta[4][0][34]  = A[4][0][34] ^ D[4][34];
    assign A_theta[4][0][35]  = A[4][0][35] ^ D[4][35];
    assign A_theta[4][0][36]  = A[4][0][36] ^ D[4][36];
    assign A_theta[4][0][37]  = A[4][0][37] ^ D[4][37];
    assign A_theta[4][0][38]  = A[4][0][38] ^ D[4][38];
    assign A_theta[4][0][39]  = A[4][0][39] ^ D[4][39];
    assign A_theta[4][0][40]  = A[4][0][40] ^ D[4][40];
    assign A_theta[4][0][41]  = A[4][0][41] ^ D[4][41];
    assign A_theta[4][0][42]  = A[4][0][42] ^ D[4][42];
    assign A_theta[4][0][43]  = A[4][0][43] ^ D[4][43];
    assign A_theta[4][0][44]  = A[4][0][44] ^ D[4][44];
    assign A_theta[4][0][45]  = A[4][0][45] ^ D[4][45];
    assign A_theta[4][0][46]  = A[4][0][46] ^ D[4][46];
    assign A_theta[4][0][47]  = A[4][0][47] ^ D[4][47];
    assign A_theta[4][0][48]  = A[4][0][48] ^ D[4][48];
    assign A_theta[4][0][49]  = A[4][0][49] ^ D[4][49];
    assign A_theta[4][0][50]  = A[4][0][50] ^ D[4][50];
    assign A_theta[4][0][51]  = A[4][0][51] ^ D[4][51];
    assign A_theta[4][0][52]  = A[4][0][52] ^ D[4][52];
    assign A_theta[4][0][53]  = A[4][0][53] ^ D[4][53];
    assign A_theta[4][0][54]  = A[4][0][54] ^ D[4][54];
    assign A_theta[4][0][55]  = A[4][0][55] ^ D[4][55];
    assign A_theta[4][0][56]  = A[4][0][56] ^ D[4][56];
    assign A_theta[4][0][57]  = A[4][0][57] ^ D[4][57];
    assign A_theta[4][0][58]  = A[4][0][58] ^ D[4][58];
    assign A_theta[4][0][59]  = A[4][0][59] ^ D[4][59];
    assign A_theta[4][0][60]  = A[4][0][60] ^ D[4][60];
    assign A_theta[4][0][61]  = A[4][0][61] ^ D[4][61];
    assign A_theta[4][0][62]  = A[4][0][62] ^ D[4][62];
    assign A_theta[4][0][63]  = A[4][0][63] ^ D[4][63];
    assign A_theta[4][1][0]  = A[4][1][0] ^ D[4][0];
    assign A_theta[4][1][1]  = A[4][1][1] ^ D[4][1];
    assign A_theta[4][1][2]  = A[4][1][2] ^ D[4][2];
    assign A_theta[4][1][3]  = A[4][1][3] ^ D[4][3];
    assign A_theta[4][1][4]  = A[4][1][4] ^ D[4][4];
    assign A_theta[4][1][5]  = A[4][1][5] ^ D[4][5];
    assign A_theta[4][1][6]  = A[4][1][6] ^ D[4][6];
    assign A_theta[4][1][7]  = A[4][1][7] ^ D[4][7];
    assign A_theta[4][1][8]  = A[4][1][8] ^ D[4][8];
    assign A_theta[4][1][9]  = A[4][1][9] ^ D[4][9];
    assign A_theta[4][1][10]  = A[4][1][10] ^ D[4][10];
    assign A_theta[4][1][11]  = A[4][1][11] ^ D[4][11];
    assign A_theta[4][1][12]  = A[4][1][12] ^ D[4][12];
    assign A_theta[4][1][13]  = A[4][1][13] ^ D[4][13];
    assign A_theta[4][1][14]  = A[4][1][14] ^ D[4][14];
    assign A_theta[4][1][15]  = A[4][1][15] ^ D[4][15];
    assign A_theta[4][1][16]  = A[4][1][16] ^ D[4][16];
    assign A_theta[4][1][17]  = A[4][1][17] ^ D[4][17];
    assign A_theta[4][1][18]  = A[4][1][18] ^ D[4][18];
    assign A_theta[4][1][19]  = A[4][1][19] ^ D[4][19];
    assign A_theta[4][1][20]  = A[4][1][20] ^ D[4][20];
    assign A_theta[4][1][21]  = A[4][1][21] ^ D[4][21];
    assign A_theta[4][1][22]  = A[4][1][22] ^ D[4][22];
    assign A_theta[4][1][23]  = A[4][1][23] ^ D[4][23];
    assign A_theta[4][1][24]  = A[4][1][24] ^ D[4][24];
    assign A_theta[4][1][25]  = A[4][1][25] ^ D[4][25];
    assign A_theta[4][1][26]  = A[4][1][26] ^ D[4][26];
    assign A_theta[4][1][27]  = A[4][1][27] ^ D[4][27];
    assign A_theta[4][1][28]  = A[4][1][28] ^ D[4][28];
    assign A_theta[4][1][29]  = A[4][1][29] ^ D[4][29];
    assign A_theta[4][1][30]  = A[4][1][30] ^ D[4][30];
    assign A_theta[4][1][31]  = A[4][1][31] ^ D[4][31];
    assign A_theta[4][1][32]  = A[4][1][32] ^ D[4][32];
    assign A_theta[4][1][33]  = A[4][1][33] ^ D[4][33];
    assign A_theta[4][1][34]  = A[4][1][34] ^ D[4][34];
    assign A_theta[4][1][35]  = A[4][1][35] ^ D[4][35];
    assign A_theta[4][1][36]  = A[4][1][36] ^ D[4][36];
    assign A_theta[4][1][37]  = A[4][1][37] ^ D[4][37];
    assign A_theta[4][1][38]  = A[4][1][38] ^ D[4][38];
    assign A_theta[4][1][39]  = A[4][1][39] ^ D[4][39];
    assign A_theta[4][1][40]  = A[4][1][40] ^ D[4][40];
    assign A_theta[4][1][41]  = A[4][1][41] ^ D[4][41];
    assign A_theta[4][1][42]  = A[4][1][42] ^ D[4][42];
    assign A_theta[4][1][43]  = A[4][1][43] ^ D[4][43];
    assign A_theta[4][1][44]  = A[4][1][44] ^ D[4][44];
    assign A_theta[4][1][45]  = A[4][1][45] ^ D[4][45];
    assign A_theta[4][1][46]  = A[4][1][46] ^ D[4][46];
    assign A_theta[4][1][47]  = A[4][1][47] ^ D[4][47];
    assign A_theta[4][1][48]  = A[4][1][48] ^ D[4][48];
    assign A_theta[4][1][49]  = A[4][1][49] ^ D[4][49];
    assign A_theta[4][1][50]  = A[4][1][50] ^ D[4][50];
    assign A_theta[4][1][51]  = A[4][1][51] ^ D[4][51];
    assign A_theta[4][1][52]  = A[4][1][52] ^ D[4][52];
    assign A_theta[4][1][53]  = A[4][1][53] ^ D[4][53];
    assign A_theta[4][1][54]  = A[4][1][54] ^ D[4][54];
    assign A_theta[4][1][55]  = A[4][1][55] ^ D[4][55];
    assign A_theta[4][1][56]  = A[4][1][56] ^ D[4][56];
    assign A_theta[4][1][57]  = A[4][1][57] ^ D[4][57];
    assign A_theta[4][1][58]  = A[4][1][58] ^ D[4][58];
    assign A_theta[4][1][59]  = A[4][1][59] ^ D[4][59];
    assign A_theta[4][1][60]  = A[4][1][60] ^ D[4][60];
    assign A_theta[4][1][61]  = A[4][1][61] ^ D[4][61];
    assign A_theta[4][1][62]  = A[4][1][62] ^ D[4][62];
    assign A_theta[4][1][63]  = A[4][1][63] ^ D[4][63];
    assign A_theta[4][2][0]  = A[4][2][0] ^ D[4][0];
    assign A_theta[4][2][1]  = A[4][2][1] ^ D[4][1];
    assign A_theta[4][2][2]  = A[4][2][2] ^ D[4][2];
    assign A_theta[4][2][3]  = A[4][2][3] ^ D[4][3];
    assign A_theta[4][2][4]  = A[4][2][4] ^ D[4][4];
    assign A_theta[4][2][5]  = A[4][2][5] ^ D[4][5];
    assign A_theta[4][2][6]  = A[4][2][6] ^ D[4][6];
    assign A_theta[4][2][7]  = A[4][2][7] ^ D[4][7];
    assign A_theta[4][2][8]  = A[4][2][8] ^ D[4][8];
    assign A_theta[4][2][9]  = A[4][2][9] ^ D[4][9];
    assign A_theta[4][2][10]  = A[4][2][10] ^ D[4][10];
    assign A_theta[4][2][11]  = A[4][2][11] ^ D[4][11];
    assign A_theta[4][2][12]  = A[4][2][12] ^ D[4][12];
    assign A_theta[4][2][13]  = A[4][2][13] ^ D[4][13];
    assign A_theta[4][2][14]  = A[4][2][14] ^ D[4][14];
    assign A_theta[4][2][15]  = A[4][2][15] ^ D[4][15];
    assign A_theta[4][2][16]  = A[4][2][16] ^ D[4][16];
    assign A_theta[4][2][17]  = A[4][2][17] ^ D[4][17];
    assign A_theta[4][2][18]  = A[4][2][18] ^ D[4][18];
    assign A_theta[4][2][19]  = A[4][2][19] ^ D[4][19];
    assign A_theta[4][2][20]  = A[4][2][20] ^ D[4][20];
    assign A_theta[4][2][21]  = A[4][2][21] ^ D[4][21];
    assign A_theta[4][2][22]  = A[4][2][22] ^ D[4][22];
    assign A_theta[4][2][23]  = A[4][2][23] ^ D[4][23];
    assign A_theta[4][2][24]  = A[4][2][24] ^ D[4][24];
    assign A_theta[4][2][25]  = A[4][2][25] ^ D[4][25];
    assign A_theta[4][2][26]  = A[4][2][26] ^ D[4][26];
    assign A_theta[4][2][27]  = A[4][2][27] ^ D[4][27];
    assign A_theta[4][2][28]  = A[4][2][28] ^ D[4][28];
    assign A_theta[4][2][29]  = A[4][2][29] ^ D[4][29];
    assign A_theta[4][2][30]  = A[4][2][30] ^ D[4][30];
    assign A_theta[4][2][31]  = A[4][2][31] ^ D[4][31];
    assign A_theta[4][2][32]  = A[4][2][32] ^ D[4][32];
    assign A_theta[4][2][33]  = A[4][2][33] ^ D[4][33];
    assign A_theta[4][2][34]  = A[4][2][34] ^ D[4][34];
    assign A_theta[4][2][35]  = A[4][2][35] ^ D[4][35];
    assign A_theta[4][2][36]  = A[4][2][36] ^ D[4][36];
    assign A_theta[4][2][37]  = A[4][2][37] ^ D[4][37];
    assign A_theta[4][2][38]  = A[4][2][38] ^ D[4][38];
    assign A_theta[4][2][39]  = A[4][2][39] ^ D[4][39];
    assign A_theta[4][2][40]  = A[4][2][40] ^ D[4][40];
    assign A_theta[4][2][41]  = A[4][2][41] ^ D[4][41];
    assign A_theta[4][2][42]  = A[4][2][42] ^ D[4][42];
    assign A_theta[4][2][43]  = A[4][2][43] ^ D[4][43];
    assign A_theta[4][2][44]  = A[4][2][44] ^ D[4][44];
    assign A_theta[4][2][45]  = A[4][2][45] ^ D[4][45];
    assign A_theta[4][2][46]  = A[4][2][46] ^ D[4][46];
    assign A_theta[4][2][47]  = A[4][2][47] ^ D[4][47];
    assign A_theta[4][2][48]  = A[4][2][48] ^ D[4][48];
    assign A_theta[4][2][49]  = A[4][2][49] ^ D[4][49];
    assign A_theta[4][2][50]  = A[4][2][50] ^ D[4][50];
    assign A_theta[4][2][51]  = A[4][2][51] ^ D[4][51];
    assign A_theta[4][2][52]  = A[4][2][52] ^ D[4][52];
    assign A_theta[4][2][53]  = A[4][2][53] ^ D[4][53];
    assign A_theta[4][2][54]  = A[4][2][54] ^ D[4][54];
    assign A_theta[4][2][55]  = A[4][2][55] ^ D[4][55];
    assign A_theta[4][2][56]  = A[4][2][56] ^ D[4][56];
    assign A_theta[4][2][57]  = A[4][2][57] ^ D[4][57];
    assign A_theta[4][2][58]  = A[4][2][58] ^ D[4][58];
    assign A_theta[4][2][59]  = A[4][2][59] ^ D[4][59];
    assign A_theta[4][2][60]  = A[4][2][60] ^ D[4][60];
    assign A_theta[4][2][61]  = A[4][2][61] ^ D[4][61];
    assign A_theta[4][2][62]  = A[4][2][62] ^ D[4][62];
    assign A_theta[4][2][63]  = A[4][2][63] ^ D[4][63];
    assign A_theta[4][3][0]  = A[4][3][0] ^ D[4][0];
    assign A_theta[4][3][1]  = A[4][3][1] ^ D[4][1];
    assign A_theta[4][3][2]  = A[4][3][2] ^ D[4][2];
    assign A_theta[4][3][3]  = A[4][3][3] ^ D[4][3];
    assign A_theta[4][3][4]  = A[4][3][4] ^ D[4][4];
    assign A_theta[4][3][5]  = A[4][3][5] ^ D[4][5];
    assign A_theta[4][3][6]  = A[4][3][6] ^ D[4][6];
    assign A_theta[4][3][7]  = A[4][3][7] ^ D[4][7];
    assign A_theta[4][3][8]  = A[4][3][8] ^ D[4][8];
    assign A_theta[4][3][9]  = A[4][3][9] ^ D[4][9];
    assign A_theta[4][3][10]  = A[4][3][10] ^ D[4][10];
    assign A_theta[4][3][11]  = A[4][3][11] ^ D[4][11];
    assign A_theta[4][3][12]  = A[4][3][12] ^ D[4][12];
    assign A_theta[4][3][13]  = A[4][3][13] ^ D[4][13];
    assign A_theta[4][3][14]  = A[4][3][14] ^ D[4][14];
    assign A_theta[4][3][15]  = A[4][3][15] ^ D[4][15];
    assign A_theta[4][3][16]  = A[4][3][16] ^ D[4][16];
    assign A_theta[4][3][17]  = A[4][3][17] ^ D[4][17];
    assign A_theta[4][3][18]  = A[4][3][18] ^ D[4][18];
    assign A_theta[4][3][19]  = A[4][3][19] ^ D[4][19];
    assign A_theta[4][3][20]  = A[4][3][20] ^ D[4][20];
    assign A_theta[4][3][21]  = A[4][3][21] ^ D[4][21];
    assign A_theta[4][3][22]  = A[4][3][22] ^ D[4][22];
    assign A_theta[4][3][23]  = A[4][3][23] ^ D[4][23];
    assign A_theta[4][3][24]  = A[4][3][24] ^ D[4][24];
    assign A_theta[4][3][25]  = A[4][3][25] ^ D[4][25];
    assign A_theta[4][3][26]  = A[4][3][26] ^ D[4][26];
    assign A_theta[4][3][27]  = A[4][3][27] ^ D[4][27];
    assign A_theta[4][3][28]  = A[4][3][28] ^ D[4][28];
    assign A_theta[4][3][29]  = A[4][3][29] ^ D[4][29];
    assign A_theta[4][3][30]  = A[4][3][30] ^ D[4][30];
    assign A_theta[4][3][31]  = A[4][3][31] ^ D[4][31];
    assign A_theta[4][3][32]  = A[4][3][32] ^ D[4][32];
    assign A_theta[4][3][33]  = A[4][3][33] ^ D[4][33];
    assign A_theta[4][3][34]  = A[4][3][34] ^ D[4][34];
    assign A_theta[4][3][35]  = A[4][3][35] ^ D[4][35];
    assign A_theta[4][3][36]  = A[4][3][36] ^ D[4][36];
    assign A_theta[4][3][37]  = A[4][3][37] ^ D[4][37];
    assign A_theta[4][3][38]  = A[4][3][38] ^ D[4][38];
    assign A_theta[4][3][39]  = A[4][3][39] ^ D[4][39];
    assign A_theta[4][3][40]  = A[4][3][40] ^ D[4][40];
    assign A_theta[4][3][41]  = A[4][3][41] ^ D[4][41];
    assign A_theta[4][3][42]  = A[4][3][42] ^ D[4][42];
    assign A_theta[4][3][43]  = A[4][3][43] ^ D[4][43];
    assign A_theta[4][3][44]  = A[4][3][44] ^ D[4][44];
    assign A_theta[4][3][45]  = A[4][3][45] ^ D[4][45];
    assign A_theta[4][3][46]  = A[4][3][46] ^ D[4][46];
    assign A_theta[4][3][47]  = A[4][3][47] ^ D[4][47];
    assign A_theta[4][3][48]  = A[4][3][48] ^ D[4][48];
    assign A_theta[4][3][49]  = A[4][3][49] ^ D[4][49];
    assign A_theta[4][3][50]  = A[4][3][50] ^ D[4][50];
    assign A_theta[4][3][51]  = A[4][3][51] ^ D[4][51];
    assign A_theta[4][3][52]  = A[4][3][52] ^ D[4][52];
    assign A_theta[4][3][53]  = A[4][3][53] ^ D[4][53];
    assign A_theta[4][3][54]  = A[4][3][54] ^ D[4][54];
    assign A_theta[4][3][55]  = A[4][3][55] ^ D[4][55];
    assign A_theta[4][3][56]  = A[4][3][56] ^ D[4][56];
    assign A_theta[4][3][57]  = A[4][3][57] ^ D[4][57];
    assign A_theta[4][3][58]  = A[4][3][58] ^ D[4][58];
    assign A_theta[4][3][59]  = A[4][3][59] ^ D[4][59];
    assign A_theta[4][3][60]  = A[4][3][60] ^ D[4][60];
    assign A_theta[4][3][61]  = A[4][3][61] ^ D[4][61];
    assign A_theta[4][3][62]  = A[4][3][62] ^ D[4][62];
    assign A_theta[4][3][63]  = A[4][3][63] ^ D[4][63];
    assign A_theta[4][4][0]  = A[4][4][0] ^ D[4][0];
    assign A_theta[4][4][1]  = A[4][4][1] ^ D[4][1];
    assign A_theta[4][4][2]  = A[4][4][2] ^ D[4][2];
    assign A_theta[4][4][3]  = A[4][4][3] ^ D[4][3];
    assign A_theta[4][4][4]  = A[4][4][4] ^ D[4][4];
    assign A_theta[4][4][5]  = A[4][4][5] ^ D[4][5];
    assign A_theta[4][4][6]  = A[4][4][6] ^ D[4][6];
    assign A_theta[4][4][7]  = A[4][4][7] ^ D[4][7];
    assign A_theta[4][4][8]  = A[4][4][8] ^ D[4][8];
    assign A_theta[4][4][9]  = A[4][4][9] ^ D[4][9];
    assign A_theta[4][4][10]  = A[4][4][10] ^ D[4][10];
    assign A_theta[4][4][11]  = A[4][4][11] ^ D[4][11];
    assign A_theta[4][4][12]  = A[4][4][12] ^ D[4][12];
    assign A_theta[4][4][13]  = A[4][4][13] ^ D[4][13];
    assign A_theta[4][4][14]  = A[4][4][14] ^ D[4][14];
    assign A_theta[4][4][15]  = A[4][4][15] ^ D[4][15];
    assign A_theta[4][4][16]  = A[4][4][16] ^ D[4][16];
    assign A_theta[4][4][17]  = A[4][4][17] ^ D[4][17];
    assign A_theta[4][4][18]  = A[4][4][18] ^ D[4][18];
    assign A_theta[4][4][19]  = A[4][4][19] ^ D[4][19];
    assign A_theta[4][4][20]  = A[4][4][20] ^ D[4][20];
    assign A_theta[4][4][21]  = A[4][4][21] ^ D[4][21];
    assign A_theta[4][4][22]  = A[4][4][22] ^ D[4][22];
    assign A_theta[4][4][23]  = A[4][4][23] ^ D[4][23];
    assign A_theta[4][4][24]  = A[4][4][24] ^ D[4][24];
    assign A_theta[4][4][25]  = A[4][4][25] ^ D[4][25];
    assign A_theta[4][4][26]  = A[4][4][26] ^ D[4][26];
    assign A_theta[4][4][27]  = A[4][4][27] ^ D[4][27];
    assign A_theta[4][4][28]  = A[4][4][28] ^ D[4][28];
    assign A_theta[4][4][29]  = A[4][4][29] ^ D[4][29];
    assign A_theta[4][4][30]  = A[4][4][30] ^ D[4][30];
    assign A_theta[4][4][31]  = A[4][4][31] ^ D[4][31];
    assign A_theta[4][4][32]  = A[4][4][32] ^ D[4][32];
    assign A_theta[4][4][33]  = A[4][4][33] ^ D[4][33];
    assign A_theta[4][4][34]  = A[4][4][34] ^ D[4][34];
    assign A_theta[4][4][35]  = A[4][4][35] ^ D[4][35];
    assign A_theta[4][4][36]  = A[4][4][36] ^ D[4][36];
    assign A_theta[4][4][37]  = A[4][4][37] ^ D[4][37];
    assign A_theta[4][4][38]  = A[4][4][38] ^ D[4][38];
    assign A_theta[4][4][39]  = A[4][4][39] ^ D[4][39];
    assign A_theta[4][4][40]  = A[4][4][40] ^ D[4][40];
    assign A_theta[4][4][41]  = A[4][4][41] ^ D[4][41];
    assign A_theta[4][4][42]  = A[4][4][42] ^ D[4][42];
    assign A_theta[4][4][43]  = A[4][4][43] ^ D[4][43];
    assign A_theta[4][4][44]  = A[4][4][44] ^ D[4][44];
    assign A_theta[4][4][45]  = A[4][4][45] ^ D[4][45];
    assign A_theta[4][4][46]  = A[4][4][46] ^ D[4][46];
    assign A_theta[4][4][47]  = A[4][4][47] ^ D[4][47];
    assign A_theta[4][4][48]  = A[4][4][48] ^ D[4][48];
    assign A_theta[4][4][49]  = A[4][4][49] ^ D[4][49];
    assign A_theta[4][4][50]  = A[4][4][50] ^ D[4][50];
    assign A_theta[4][4][51]  = A[4][4][51] ^ D[4][51];
    assign A_theta[4][4][52]  = A[4][4][52] ^ D[4][52];
    assign A_theta[4][4][53]  = A[4][4][53] ^ D[4][53];
    assign A_theta[4][4][54]  = A[4][4][54] ^ D[4][54];
    assign A_theta[4][4][55]  = A[4][4][55] ^ D[4][55];
    assign A_theta[4][4][56]  = A[4][4][56] ^ D[4][56];
    assign A_theta[4][4][57]  = A[4][4][57] ^ D[4][57];
    assign A_theta[4][4][58]  = A[4][4][58] ^ D[4][58];
    assign A_theta[4][4][59]  = A[4][4][59] ^ D[4][59];
    assign A_theta[4][4][60]  = A[4][4][60] ^ D[4][60];
    assign A_theta[4][4][61]  = A[4][4][61] ^ D[4][61];
    assign A_theta[4][4][62]  = A[4][4][62] ^ D[4][62];
    assign A_theta[4][4][63]  = A[4][4][63] ^ D[4][63];
//--------------------------- RHO ---------------------------
    // Step 1: Copy A[0][0][z] to A_rho[0][0][z]
    assign A_rho[0][0][0]    = A[0][0][0];
    assign A_rho[0][0][1]    = A[0][0][1];
    assign A_rho[0][0][2]    = A[0][0][2];
    assign A_rho[0][0][3]    = A[0][0][3];
    assign A_rho[0][0][4]    = A[0][0][4];
    assign A_rho[0][0][5]    = A[0][0][5];
    assign A_rho[0][0][6]    = A[0][0][6];
    assign A_rho[0][0][7]    = A[0][0][7];
    assign A_rho[0][0][8]    = A[0][0][8];
    assign A_rho[0][0][9]    = A[0][0][9];
    assign A_rho[0][0][10]    = A[0][0][10];
    assign A_rho[0][0][11]    = A[0][0][11];
    assign A_rho[0][0][12]    = A[0][0][12];
    assign A_rho[0][0][13]    = A[0][0][13];
    assign A_rho[0][0][14]    = A[0][0][14];
    assign A_rho[0][0][15]    = A[0][0][15];
    assign A_rho[0][0][16]    = A[0][0][16];
    assign A_rho[0][0][17]    = A[0][0][17];
    assign A_rho[0][0][18]    = A[0][0][18];
    assign A_rho[0][0][19]    = A[0][0][19];
    assign A_rho[0][0][20]    = A[0][0][20];
    assign A_rho[0][0][21]    = A[0][0][21];
    assign A_rho[0][0][22]    = A[0][0][22];
    assign A_rho[0][0][23]    = A[0][0][23];
    assign A_rho[0][0][24]    = A[0][0][24];
    assign A_rho[0][0][25]    = A[0][0][25];
    assign A_rho[0][0][26]    = A[0][0][26];
    assign A_rho[0][0][27]    = A[0][0][27];
    assign A_rho[0][0][28]    = A[0][0][28];
    assign A_rho[0][0][29]    = A[0][0][29];
    assign A_rho[0][0][30]    = A[0][0][30];
    assign A_rho[0][0][31]    = A[0][0][31];
    assign A_rho[0][0][32]    = A[0][0][32];
    assign A_rho[0][0][33]    = A[0][0][33];
    assign A_rho[0][0][34]    = A[0][0][34];
    assign A_rho[0][0][35]    = A[0][0][35];
    assign A_rho[0][0][36]    = A[0][0][36];
    assign A_rho[0][0][37]    = A[0][0][37];
    assign A_rho[0][0][38]    = A[0][0][38];
    assign A_rho[0][0][39]    = A[0][0][39];
    assign A_rho[0][0][40]    = A[0][0][40];
    assign A_rho[0][0][41]    = A[0][0][41];
    assign A_rho[0][0][42]    = A[0][0][42];
    assign A_rho[0][0][43]    = A[0][0][43];
    assign A_rho[0][0][44]    = A[0][0][44];
    assign A_rho[0][0][45]    = A[0][0][45];
    assign A_rho[0][0][46]    = A[0][0][46];
    assign A_rho[0][0][47]    = A[0][0][47];
    assign A_rho[0][0][48]    = A[0][0][48];
    assign A_rho[0][0][49]    = A[0][0][49];
    assign A_rho[0][0][50]    = A[0][0][50];
    assign A_rho[0][0][51]    = A[0][0][51];
    assign A_rho[0][0][52]    = A[0][0][52];
    assign A_rho[0][0][53]    = A[0][0][53];
    assign A_rho[0][0][54]    = A[0][0][54];
    assign A_rho[0][0][55]    = A[0][0][55];
    assign A_rho[0][0][56]    = A[0][0][56];
    assign A_rho[0][0][57]    = A[0][0][57];
    assign A_rho[0][0][58]    = A[0][0][58];
    assign A_rho[0][0][59]    = A[0][0][59];
    assign A_rho[0][0][60]    = A[0][0][60];
    assign A_rho[0][0][61]    = A[0][0][61];
    assign A_rho[0][0][62]    = A[0][0][62];
    assign A_rho[0][0][63]    = A[0][0][63];

    // Step 2: Transformations for other lanes
    assign A_rho[1][0][0]    = A[1][0][63];
    assign A_rho[1][0][1]    = A[1][0][0];
    assign A_rho[1][0][2]    = A[1][0][1];
    assign A_rho[1][0][3]    = A[1][0][2];
    assign A_rho[1][0][4]    = A[1][0][3];
    assign A_rho[1][0][5]    = A[1][0][4];
    assign A_rho[1][0][6]    = A[1][0][5];
    assign A_rho[1][0][7]    = A[1][0][6];
    assign A_rho[1][0][8]    = A[1][0][7];
    assign A_rho[1][0][9]    = A[1][0][8];
    assign A_rho[1][0][10]    = A[1][0][9];
    assign A_rho[1][0][11]    = A[1][0][10];
    assign A_rho[1][0][12]    = A[1][0][11];
    assign A_rho[1][0][13]    = A[1][0][12];
    assign A_rho[1][0][14]    = A[1][0][13];
    assign A_rho[1][0][15]    = A[1][0][14];
    assign A_rho[1][0][16]    = A[1][0][15];
    assign A_rho[1][0][17]    = A[1][0][16];
    assign A_rho[1][0][18]    = A[1][0][17];
    assign A_rho[1][0][19]    = A[1][0][18];
    assign A_rho[1][0][20]    = A[1][0][19];
    assign A_rho[1][0][21]    = A[1][0][20];
    assign A_rho[1][0][22]    = A[1][0][21];
    assign A_rho[1][0][23]    = A[1][0][22];
    assign A_rho[1][0][24]    = A[1][0][23];
    assign A_rho[1][0][25]    = A[1][0][24];
    assign A_rho[1][0][26]    = A[1][0][25];
    assign A_rho[1][0][27]    = A[1][0][26];
    assign A_rho[1][0][28]    = A[1][0][27];
    assign A_rho[1][0][29]    = A[1][0][28];
    assign A_rho[1][0][30]    = A[1][0][29];
    assign A_rho[1][0][31]    = A[1][0][30];
    assign A_rho[1][0][32]    = A[1][0][31];
    assign A_rho[1][0][33]    = A[1][0][32];
    assign A_rho[1][0][34]    = A[1][0][33];
    assign A_rho[1][0][35]    = A[1][0][34];
    assign A_rho[1][0][36]    = A[1][0][35];
    assign A_rho[1][0][37]    = A[1][0][36];
    assign A_rho[1][0][38]    = A[1][0][37];
    assign A_rho[1][0][39]    = A[1][0][38];
    assign A_rho[1][0][40]    = A[1][0][39];
    assign A_rho[1][0][41]    = A[1][0][40];
    assign A_rho[1][0][42]    = A[1][0][41];
    assign A_rho[1][0][43]    = A[1][0][42];
    assign A_rho[1][0][44]    = A[1][0][43];
    assign A_rho[1][0][45]    = A[1][0][44];
    assign A_rho[1][0][46]    = A[1][0][45];
    assign A_rho[1][0][47]    = A[1][0][46];
    assign A_rho[1][0][48]    = A[1][0][47];
    assign A_rho[1][0][49]    = A[1][0][48];
    assign A_rho[1][0][50]    = A[1][0][49];
    assign A_rho[1][0][51]    = A[1][0][50];
    assign A_rho[1][0][52]    = A[1][0][51];
    assign A_rho[1][0][53]    = A[1][0][52];
    assign A_rho[1][0][54]    = A[1][0][53];
    assign A_rho[1][0][55]    = A[1][0][54];
    assign A_rho[1][0][56]    = A[1][0][55];
    assign A_rho[1][0][57]    = A[1][0][56];
    assign A_rho[1][0][58]    = A[1][0][57];
    assign A_rho[1][0][59]    = A[1][0][58];
    assign A_rho[1][0][60]    = A[1][0][59];
    assign A_rho[1][0][61]    = A[1][0][60];
    assign A_rho[1][0][62]    = A[1][0][61];
    assign A_rho[1][0][63]    = A[1][0][62];
    assign A_rho[0][2][0]    = A[0][2][61];
    assign A_rho[0][2][1]    = A[0][2][62];
    assign A_rho[0][2][2]    = A[0][2][63];
    assign A_rho[0][2][3]    = A[0][2][0];
    assign A_rho[0][2][4]    = A[0][2][1];
    assign A_rho[0][2][5]    = A[0][2][2];
    assign A_rho[0][2][6]    = A[0][2][3];
    assign A_rho[0][2][7]    = A[0][2][4];
    assign A_rho[0][2][8]    = A[0][2][5];
    assign A_rho[0][2][9]    = A[0][2][6];
    assign A_rho[0][2][10]    = A[0][2][7];
    assign A_rho[0][2][11]    = A[0][2][8];
    assign A_rho[0][2][12]    = A[0][2][9];
    assign A_rho[0][2][13]    = A[0][2][10];
    assign A_rho[0][2][14]    = A[0][2][11];
    assign A_rho[0][2][15]    = A[0][2][12];
    assign A_rho[0][2][16]    = A[0][2][13];
    assign A_rho[0][2][17]    = A[0][2][14];
    assign A_rho[0][2][18]    = A[0][2][15];
    assign A_rho[0][2][19]    = A[0][2][16];
    assign A_rho[0][2][20]    = A[0][2][17];
    assign A_rho[0][2][21]    = A[0][2][18];
    assign A_rho[0][2][22]    = A[0][2][19];
    assign A_rho[0][2][23]    = A[0][2][20];
    assign A_rho[0][2][24]    = A[0][2][21];
    assign A_rho[0][2][25]    = A[0][2][22];
    assign A_rho[0][2][26]    = A[0][2][23];
    assign A_rho[0][2][27]    = A[0][2][24];
    assign A_rho[0][2][28]    = A[0][2][25];
    assign A_rho[0][2][29]    = A[0][2][26];
    assign A_rho[0][2][30]    = A[0][2][27];
    assign A_rho[0][2][31]    = A[0][2][28];
    assign A_rho[0][2][32]    = A[0][2][29];
    assign A_rho[0][2][33]    = A[0][2][30];
    assign A_rho[0][2][34]    = A[0][2][31];
    assign A_rho[0][2][35]    = A[0][2][32];
    assign A_rho[0][2][36]    = A[0][2][33];
    assign A_rho[0][2][37]    = A[0][2][34];
    assign A_rho[0][2][38]    = A[0][2][35];
    assign A_rho[0][2][39]    = A[0][2][36];
    assign A_rho[0][2][40]    = A[0][2][37];
    assign A_rho[0][2][41]    = A[0][2][38];
    assign A_rho[0][2][42]    = A[0][2][39];
    assign A_rho[0][2][43]    = A[0][2][40];
    assign A_rho[0][2][44]    = A[0][2][41];
    assign A_rho[0][2][45]    = A[0][2][42];
    assign A_rho[0][2][46]    = A[0][2][43];
    assign A_rho[0][2][47]    = A[0][2][44];
    assign A_rho[0][2][48]    = A[0][2][45];
    assign A_rho[0][2][49]    = A[0][2][46];
    assign A_rho[0][2][50]    = A[0][2][47];
    assign A_rho[0][2][51]    = A[0][2][48];
    assign A_rho[0][2][52]    = A[0][2][49];
    assign A_rho[0][2][53]    = A[0][2][50];
    assign A_rho[0][2][54]    = A[0][2][51];
    assign A_rho[0][2][55]    = A[0][2][52];
    assign A_rho[0][2][56]    = A[0][2][53];
    assign A_rho[0][2][57]    = A[0][2][54];
    assign A_rho[0][2][58]    = A[0][2][55];
    assign A_rho[0][2][59]    = A[0][2][56];
    assign A_rho[0][2][60]    = A[0][2][57];
    assign A_rho[0][2][61]    = A[0][2][58];
    assign A_rho[0][2][62]    = A[0][2][59];
    assign A_rho[0][2][63]    = A[0][2][60];
    assign A_rho[2][1][0]    = A[2][1][58];
    assign A_rho[2][1][1]    = A[2][1][59];
    assign A_rho[2][1][2]    = A[2][1][60];
    assign A_rho[2][1][3]    = A[2][1][61];
    assign A_rho[2][1][4]    = A[2][1][62];
    assign A_rho[2][1][5]    = A[2][1][63];
    assign A_rho[2][1][6]    = A[2][1][0];
    assign A_rho[2][1][7]    = A[2][1][1];
    assign A_rho[2][1][8]    = A[2][1][2];
    assign A_rho[2][1][9]    = A[2][1][3];
    assign A_rho[2][1][10]    = A[2][1][4];
    assign A_rho[2][1][11]    = A[2][1][5];
    assign A_rho[2][1][12]    = A[2][1][6];
    assign A_rho[2][1][13]    = A[2][1][7];
    assign A_rho[2][1][14]    = A[2][1][8];
    assign A_rho[2][1][15]    = A[2][1][9];
    assign A_rho[2][1][16]    = A[2][1][10];
    assign A_rho[2][1][17]    = A[2][1][11];
    assign A_rho[2][1][18]    = A[2][1][12];
    assign A_rho[2][1][19]    = A[2][1][13];
    assign A_rho[2][1][20]    = A[2][1][14];
    assign A_rho[2][1][21]    = A[2][1][15];
    assign A_rho[2][1][22]    = A[2][1][16];
    assign A_rho[2][1][23]    = A[2][1][17];
    assign A_rho[2][1][24]    = A[2][1][18];
    assign A_rho[2][1][25]    = A[2][1][19];
    assign A_rho[2][1][26]    = A[2][1][20];
    assign A_rho[2][1][27]    = A[2][1][21];
    assign A_rho[2][1][28]    = A[2][1][22];
    assign A_rho[2][1][29]    = A[2][1][23];
    assign A_rho[2][1][30]    = A[2][1][24];
    assign A_rho[2][1][31]    = A[2][1][25];
    assign A_rho[2][1][32]    = A[2][1][26];
    assign A_rho[2][1][33]    = A[2][1][27];
    assign A_rho[2][1][34]    = A[2][1][28];
    assign A_rho[2][1][35]    = A[2][1][29];
    assign A_rho[2][1][36]    = A[2][1][30];
    assign A_rho[2][1][37]    = A[2][1][31];
    assign A_rho[2][1][38]    = A[2][1][32];
    assign A_rho[2][1][39]    = A[2][1][33];
    assign A_rho[2][1][40]    = A[2][1][34];
    assign A_rho[2][1][41]    = A[2][1][35];
    assign A_rho[2][1][42]    = A[2][1][36];
    assign A_rho[2][1][43]    = A[2][1][37];
    assign A_rho[2][1][44]    = A[2][1][38];
    assign A_rho[2][1][45]    = A[2][1][39];
    assign A_rho[2][1][46]    = A[2][1][40];
    assign A_rho[2][1][47]    = A[2][1][41];
    assign A_rho[2][1][48]    = A[2][1][42];
    assign A_rho[2][1][49]    = A[2][1][43];
    assign A_rho[2][1][50]    = A[2][1][44];
    assign A_rho[2][1][51]    = A[2][1][45];
    assign A_rho[2][1][52]    = A[2][1][46];
    assign A_rho[2][1][53]    = A[2][1][47];
    assign A_rho[2][1][54]    = A[2][1][48];
    assign A_rho[2][1][55]    = A[2][1][49];
    assign A_rho[2][1][56]    = A[2][1][50];
    assign A_rho[2][1][57]    = A[2][1][51];
    assign A_rho[2][1][58]    = A[2][1][52];
    assign A_rho[2][1][59]    = A[2][1][53];
    assign A_rho[2][1][60]    = A[2][1][54];
    assign A_rho[2][1][61]    = A[2][1][55];
    assign A_rho[2][1][62]    = A[2][1][56];
    assign A_rho[2][1][63]    = A[2][1][57];
    assign A_rho[1][2][0]    = A[1][2][54];
    assign A_rho[1][2][1]    = A[1][2][55];
    assign A_rho[1][2][2]    = A[1][2][56];
    assign A_rho[1][2][3]    = A[1][2][57];
    assign A_rho[1][2][4]    = A[1][2][58];
    assign A_rho[1][2][5]    = A[1][2][59];
    assign A_rho[1][2][6]    = A[1][2][60];
    assign A_rho[1][2][7]    = A[1][2][61];
    assign A_rho[1][2][8]    = A[1][2][62];
    assign A_rho[1][2][9]    = A[1][2][63];
    assign A_rho[1][2][10]    = A[1][2][0];
    assign A_rho[1][2][11]    = A[1][2][1];
    assign A_rho[1][2][12]    = A[1][2][2];
    assign A_rho[1][2][13]    = A[1][2][3];
    assign A_rho[1][2][14]    = A[1][2][4];
    assign A_rho[1][2][15]    = A[1][2][5];
    assign A_rho[1][2][16]    = A[1][2][6];
    assign A_rho[1][2][17]    = A[1][2][7];
    assign A_rho[1][2][18]    = A[1][2][8];
    assign A_rho[1][2][19]    = A[1][2][9];
    assign A_rho[1][2][20]    = A[1][2][10];
    assign A_rho[1][2][21]    = A[1][2][11];
    assign A_rho[1][2][22]    = A[1][2][12];
    assign A_rho[1][2][23]    = A[1][2][13];
    assign A_rho[1][2][24]    = A[1][2][14];
    assign A_rho[1][2][25]    = A[1][2][15];
    assign A_rho[1][2][26]    = A[1][2][16];
    assign A_rho[1][2][27]    = A[1][2][17];
    assign A_rho[1][2][28]    = A[1][2][18];
    assign A_rho[1][2][29]    = A[1][2][19];
    assign A_rho[1][2][30]    = A[1][2][20];
    assign A_rho[1][2][31]    = A[1][2][21];
    assign A_rho[1][2][32]    = A[1][2][22];
    assign A_rho[1][2][33]    = A[1][2][23];
    assign A_rho[1][2][34]    = A[1][2][24];
    assign A_rho[1][2][35]    = A[1][2][25];
    assign A_rho[1][2][36]    = A[1][2][26];
    assign A_rho[1][2][37]    = A[1][2][27];
    assign A_rho[1][2][38]    = A[1][2][28];
    assign A_rho[1][2][39]    = A[1][2][29];
    assign A_rho[1][2][40]    = A[1][2][30];
    assign A_rho[1][2][41]    = A[1][2][31];
    assign A_rho[1][2][42]    = A[1][2][32];
    assign A_rho[1][2][43]    = A[1][2][33];
    assign A_rho[1][2][44]    = A[1][2][34];
    assign A_rho[1][2][45]    = A[1][2][35];
    assign A_rho[1][2][46]    = A[1][2][36];
    assign A_rho[1][2][47]    = A[1][2][37];
    assign A_rho[1][2][48]    = A[1][2][38];
    assign A_rho[1][2][49]    = A[1][2][39];
    assign A_rho[1][2][50]    = A[1][2][40];
    assign A_rho[1][2][51]    = A[1][2][41];
    assign A_rho[1][2][52]    = A[1][2][42];
    assign A_rho[1][2][53]    = A[1][2][43];
    assign A_rho[1][2][54]    = A[1][2][44];
    assign A_rho[1][2][55]    = A[1][2][45];
    assign A_rho[1][2][56]    = A[1][2][46];
    assign A_rho[1][2][57]    = A[1][2][47];
    assign A_rho[1][2][58]    = A[1][2][48];
    assign A_rho[1][2][59]    = A[1][2][49];
    assign A_rho[1][2][60]    = A[1][2][50];
    assign A_rho[1][2][61]    = A[1][2][51];
    assign A_rho[1][2][62]    = A[1][2][52];
    assign A_rho[1][2][63]    = A[1][2][53];
    assign A_rho[2][3][0]    = A[2][3][49];
    assign A_rho[2][3][1]    = A[2][3][50];
    assign A_rho[2][3][2]    = A[2][3][51];
    assign A_rho[2][3][3]    = A[2][3][52];
    assign A_rho[2][3][4]    = A[2][3][53];
    assign A_rho[2][3][5]    = A[2][3][54];
    assign A_rho[2][3][6]    = A[2][3][55];
    assign A_rho[2][3][7]    = A[2][3][56];
    assign A_rho[2][3][8]    = A[2][3][57];
    assign A_rho[2][3][9]    = A[2][3][58];
    assign A_rho[2][3][10]    = A[2][3][59];
    assign A_rho[2][3][11]    = A[2][3][60];
    assign A_rho[2][3][12]    = A[2][3][61];
    assign A_rho[2][3][13]    = A[2][3][62];
    assign A_rho[2][3][14]    = A[2][3][63];
    assign A_rho[2][3][15]    = A[2][3][0];
    assign A_rho[2][3][16]    = A[2][3][1];
    assign A_rho[2][3][17]    = A[2][3][2];
    assign A_rho[2][3][18]    = A[2][3][3];
    assign A_rho[2][3][19]    = A[2][3][4];
    assign A_rho[2][3][20]    = A[2][3][5];
    assign A_rho[2][3][21]    = A[2][3][6];
    assign A_rho[2][3][22]    = A[2][3][7];
    assign A_rho[2][3][23]    = A[2][3][8];
    assign A_rho[2][3][24]    = A[2][3][9];
    assign A_rho[2][3][25]    = A[2][3][10];
    assign A_rho[2][3][26]    = A[2][3][11];
    assign A_rho[2][3][27]    = A[2][3][12];
    assign A_rho[2][3][28]    = A[2][3][13];
    assign A_rho[2][3][29]    = A[2][3][14];
    assign A_rho[2][3][30]    = A[2][3][15];
    assign A_rho[2][3][31]    = A[2][3][16];
    assign A_rho[2][3][32]    = A[2][3][17];
    assign A_rho[2][3][33]    = A[2][3][18];
    assign A_rho[2][3][34]    = A[2][3][19];
    assign A_rho[2][3][35]    = A[2][3][20];
    assign A_rho[2][3][36]    = A[2][3][21];
    assign A_rho[2][3][37]    = A[2][3][22];
    assign A_rho[2][3][38]    = A[2][3][23];
    assign A_rho[2][3][39]    = A[2][3][24];
    assign A_rho[2][3][40]    = A[2][3][25];
    assign A_rho[2][3][41]    = A[2][3][26];
    assign A_rho[2][3][42]    = A[2][3][27];
    assign A_rho[2][3][43]    = A[2][3][28];
    assign A_rho[2][3][44]    = A[2][3][29];
    assign A_rho[2][3][45]    = A[2][3][30];
    assign A_rho[2][3][46]    = A[2][3][31];
    assign A_rho[2][3][47]    = A[2][3][32];
    assign A_rho[2][3][48]    = A[2][3][33];
    assign A_rho[2][3][49]    = A[2][3][34];
    assign A_rho[2][3][50]    = A[2][3][35];
    assign A_rho[2][3][51]    = A[2][3][36];
    assign A_rho[2][3][52]    = A[2][3][37];
    assign A_rho[2][3][53]    = A[2][3][38];
    assign A_rho[2][3][54]    = A[2][3][39];
    assign A_rho[2][3][55]    = A[2][3][40];
    assign A_rho[2][3][56]    = A[2][3][41];
    assign A_rho[2][3][57]    = A[2][3][42];
    assign A_rho[2][3][58]    = A[2][3][43];
    assign A_rho[2][3][59]    = A[2][3][44];
    assign A_rho[2][3][60]    = A[2][3][45];
    assign A_rho[2][3][61]    = A[2][3][46];
    assign A_rho[2][3][62]    = A[2][3][47];
    assign A_rho[2][3][63]    = A[2][3][48];
    assign A_rho[3][3][0]    = A[3][3][43];
    assign A_rho[3][3][1]    = A[3][3][44];
    assign A_rho[3][3][2]    = A[3][3][45];
    assign A_rho[3][3][3]    = A[3][3][46];
    assign A_rho[3][3][4]    = A[3][3][47];
    assign A_rho[3][3][5]    = A[3][3][48];
    assign A_rho[3][3][6]    = A[3][3][49];
    assign A_rho[3][3][7]    = A[3][3][50];
    assign A_rho[3][3][8]    = A[3][3][51];
    assign A_rho[3][3][9]    = A[3][3][52];
    assign A_rho[3][3][10]    = A[3][3][53];
    assign A_rho[3][3][11]    = A[3][3][54];
    assign A_rho[3][3][12]    = A[3][3][55];
    assign A_rho[3][3][13]    = A[3][3][56];
    assign A_rho[3][3][14]    = A[3][3][57];
    assign A_rho[3][3][15]    = A[3][3][58];
    assign A_rho[3][3][16]    = A[3][3][59];
    assign A_rho[3][3][17]    = A[3][3][60];
    assign A_rho[3][3][18]    = A[3][3][61];
    assign A_rho[3][3][19]    = A[3][3][62];
    assign A_rho[3][3][20]    = A[3][3][63];
    assign A_rho[3][3][21]    = A[3][3][0];
    assign A_rho[3][3][22]    = A[3][3][1];
    assign A_rho[3][3][23]    = A[3][3][2];
    assign A_rho[3][3][24]    = A[3][3][3];
    assign A_rho[3][3][25]    = A[3][3][4];
    assign A_rho[3][3][26]    = A[3][3][5];
    assign A_rho[3][3][27]    = A[3][3][6];
    assign A_rho[3][3][28]    = A[3][3][7];
    assign A_rho[3][3][29]    = A[3][3][8];
    assign A_rho[3][3][30]    = A[3][3][9];
    assign A_rho[3][3][31]    = A[3][3][10];
    assign A_rho[3][3][32]    = A[3][3][11];
    assign A_rho[3][3][33]    = A[3][3][12];
    assign A_rho[3][3][34]    = A[3][3][13];
    assign A_rho[3][3][35]    = A[3][3][14];
    assign A_rho[3][3][36]    = A[3][3][15];
    assign A_rho[3][3][37]    = A[3][3][16];
    assign A_rho[3][3][38]    = A[3][3][17];
    assign A_rho[3][3][39]    = A[3][3][18];
    assign A_rho[3][3][40]    = A[3][3][19];
    assign A_rho[3][3][41]    = A[3][3][20];
    assign A_rho[3][3][42]    = A[3][3][21];
    assign A_rho[3][3][43]    = A[3][3][22];
    assign A_rho[3][3][44]    = A[3][3][23];
    assign A_rho[3][3][45]    = A[3][3][24];
    assign A_rho[3][3][46]    = A[3][3][25];
    assign A_rho[3][3][47]    = A[3][3][26];
    assign A_rho[3][3][48]    = A[3][3][27];
    assign A_rho[3][3][49]    = A[3][3][28];
    assign A_rho[3][3][50]    = A[3][3][29];
    assign A_rho[3][3][51]    = A[3][3][30];
    assign A_rho[3][3][52]    = A[3][3][31];
    assign A_rho[3][3][53]    = A[3][3][32];
    assign A_rho[3][3][54]    = A[3][3][33];
    assign A_rho[3][3][55]    = A[3][3][34];
    assign A_rho[3][3][56]    = A[3][3][35];
    assign A_rho[3][3][57]    = A[3][3][36];
    assign A_rho[3][3][58]    = A[3][3][37];
    assign A_rho[3][3][59]    = A[3][3][38];
    assign A_rho[3][3][60]    = A[3][3][39];
    assign A_rho[3][3][61]    = A[3][3][40];
    assign A_rho[3][3][62]    = A[3][3][41];
    assign A_rho[3][3][63]    = A[3][3][42];
    assign A_rho[3][0][0]    = A[3][0][36];
    assign A_rho[3][0][1]    = A[3][0][37];
    assign A_rho[3][0][2]    = A[3][0][38];
    assign A_rho[3][0][3]    = A[3][0][39];
    assign A_rho[3][0][4]    = A[3][0][40];
    assign A_rho[3][0][5]    = A[3][0][41];
    assign A_rho[3][0][6]    = A[3][0][42];
    assign A_rho[3][0][7]    = A[3][0][43];
    assign A_rho[3][0][8]    = A[3][0][44];
    assign A_rho[3][0][9]    = A[3][0][45];
    assign A_rho[3][0][10]    = A[3][0][46];
    assign A_rho[3][0][11]    = A[3][0][47];
    assign A_rho[3][0][12]    = A[3][0][48];
    assign A_rho[3][0][13]    = A[3][0][49];
    assign A_rho[3][0][14]    = A[3][0][50];
    assign A_rho[3][0][15]    = A[3][0][51];
    assign A_rho[3][0][16]    = A[3][0][52];
    assign A_rho[3][0][17]    = A[3][0][53];
    assign A_rho[3][0][18]    = A[3][0][54];
    assign A_rho[3][0][19]    = A[3][0][55];
    assign A_rho[3][0][20]    = A[3][0][56];
    assign A_rho[3][0][21]    = A[3][0][57];
    assign A_rho[3][0][22]    = A[3][0][58];
    assign A_rho[3][0][23]    = A[3][0][59];
    assign A_rho[3][0][24]    = A[3][0][60];
    assign A_rho[3][0][25]    = A[3][0][61];
    assign A_rho[3][0][26]    = A[3][0][62];
    assign A_rho[3][0][27]    = A[3][0][63];
    assign A_rho[3][0][28]    = A[3][0][0];
    assign A_rho[3][0][29]    = A[3][0][1];
    assign A_rho[3][0][30]    = A[3][0][2];
    assign A_rho[3][0][31]    = A[3][0][3];
    assign A_rho[3][0][32]    = A[3][0][4];
    assign A_rho[3][0][33]    = A[3][0][5];
    assign A_rho[3][0][34]    = A[3][0][6];
    assign A_rho[3][0][35]    = A[3][0][7];
    assign A_rho[3][0][36]    = A[3][0][8];
    assign A_rho[3][0][37]    = A[3][0][9];
    assign A_rho[3][0][38]    = A[3][0][10];
    assign A_rho[3][0][39]    = A[3][0][11];
    assign A_rho[3][0][40]    = A[3][0][12];
    assign A_rho[3][0][41]    = A[3][0][13];
    assign A_rho[3][0][42]    = A[3][0][14];
    assign A_rho[3][0][43]    = A[3][0][15];
    assign A_rho[3][0][44]    = A[3][0][16];
    assign A_rho[3][0][45]    = A[3][0][17];
    assign A_rho[3][0][46]    = A[3][0][18];
    assign A_rho[3][0][47]    = A[3][0][19];
    assign A_rho[3][0][48]    = A[3][0][20];
    assign A_rho[3][0][49]    = A[3][0][21];
    assign A_rho[3][0][50]    = A[3][0][22];
    assign A_rho[3][0][51]    = A[3][0][23];
    assign A_rho[3][0][52]    = A[3][0][24];
    assign A_rho[3][0][53]    = A[3][0][25];
    assign A_rho[3][0][54]    = A[3][0][26];
    assign A_rho[3][0][55]    = A[3][0][27];
    assign A_rho[3][0][56]    = A[3][0][28];
    assign A_rho[3][0][57]    = A[3][0][29];
    assign A_rho[3][0][58]    = A[3][0][30];
    assign A_rho[3][0][59]    = A[3][0][31];
    assign A_rho[3][0][60]    = A[3][0][32];
    assign A_rho[3][0][61]    = A[3][0][33];
    assign A_rho[3][0][62]    = A[3][0][34];
    assign A_rho[3][0][63]    = A[3][0][35];
    assign A_rho[0][1][0]    = A[0][1][28];
    assign A_rho[0][1][1]    = A[0][1][29];
    assign A_rho[0][1][2]    = A[0][1][30];
    assign A_rho[0][1][3]    = A[0][1][31];
    assign A_rho[0][1][4]    = A[0][1][32];
    assign A_rho[0][1][5]    = A[0][1][33];
    assign A_rho[0][1][6]    = A[0][1][34];
    assign A_rho[0][1][7]    = A[0][1][35];
    assign A_rho[0][1][8]    = A[0][1][36];
    assign A_rho[0][1][9]    = A[0][1][37];
    assign A_rho[0][1][10]    = A[0][1][38];
    assign A_rho[0][1][11]    = A[0][1][39];
    assign A_rho[0][1][12]    = A[0][1][40];
    assign A_rho[0][1][13]    = A[0][1][41];
    assign A_rho[0][1][14]    = A[0][1][42];
    assign A_rho[0][1][15]    = A[0][1][43];
    assign A_rho[0][1][16]    = A[0][1][44];
    assign A_rho[0][1][17]    = A[0][1][45];
    assign A_rho[0][1][18]    = A[0][1][46];
    assign A_rho[0][1][19]    = A[0][1][47];
    assign A_rho[0][1][20]    = A[0][1][48];
    assign A_rho[0][1][21]    = A[0][1][49];
    assign A_rho[0][1][22]    = A[0][1][50];
    assign A_rho[0][1][23]    = A[0][1][51];
    assign A_rho[0][1][24]    = A[0][1][52];
    assign A_rho[0][1][25]    = A[0][1][53];
    assign A_rho[0][1][26]    = A[0][1][54];
    assign A_rho[0][1][27]    = A[0][1][55];
    assign A_rho[0][1][28]    = A[0][1][56];
    assign A_rho[0][1][29]    = A[0][1][57];
    assign A_rho[0][1][30]    = A[0][1][58];
    assign A_rho[0][1][31]    = A[0][1][59];
    assign A_rho[0][1][32]    = A[0][1][60];
    assign A_rho[0][1][33]    = A[0][1][61];
    assign A_rho[0][1][34]    = A[0][1][62];
    assign A_rho[0][1][35]    = A[0][1][63];
    assign A_rho[0][1][36]    = A[0][1][0];
    assign A_rho[0][1][37]    = A[0][1][1];
    assign A_rho[0][1][38]    = A[0][1][2];
    assign A_rho[0][1][39]    = A[0][1][3];
    assign A_rho[0][1][40]    = A[0][1][4];
    assign A_rho[0][1][41]    = A[0][1][5];
    assign A_rho[0][1][42]    = A[0][1][6];
    assign A_rho[0][1][43]    = A[0][1][7];
    assign A_rho[0][1][44]    = A[0][1][8];
    assign A_rho[0][1][45]    = A[0][1][9];
    assign A_rho[0][1][46]    = A[0][1][10];
    assign A_rho[0][1][47]    = A[0][1][11];
    assign A_rho[0][1][48]    = A[0][1][12];
    assign A_rho[0][1][49]    = A[0][1][13];
    assign A_rho[0][1][50]    = A[0][1][14];
    assign A_rho[0][1][51]    = A[0][1][15];
    assign A_rho[0][1][52]    = A[0][1][16];
    assign A_rho[0][1][53]    = A[0][1][17];
    assign A_rho[0][1][54]    = A[0][1][18];
    assign A_rho[0][1][55]    = A[0][1][19];
    assign A_rho[0][1][56]    = A[0][1][20];
    assign A_rho[0][1][57]    = A[0][1][21];
    assign A_rho[0][1][58]    = A[0][1][22];
    assign A_rho[0][1][59]    = A[0][1][23];
    assign A_rho[0][1][60]    = A[0][1][24];
    assign A_rho[0][1][61]    = A[0][1][25];
    assign A_rho[0][1][62]    = A[0][1][26];
    assign A_rho[0][1][63]    = A[0][1][27];
    assign A_rho[1][3][0]    = A[1][3][19];
    assign A_rho[1][3][1]    = A[1][3][20];
    assign A_rho[1][3][2]    = A[1][3][21];
    assign A_rho[1][3][3]    = A[1][3][22];
    assign A_rho[1][3][4]    = A[1][3][23];
    assign A_rho[1][3][5]    = A[1][3][24];
    assign A_rho[1][3][6]    = A[1][3][25];
    assign A_rho[1][3][7]    = A[1][3][26];
    assign A_rho[1][3][8]    = A[1][3][27];
    assign A_rho[1][3][9]    = A[1][3][28];
    assign A_rho[1][3][10]    = A[1][3][29];
    assign A_rho[1][3][11]    = A[1][3][30];
    assign A_rho[1][3][12]    = A[1][3][31];
    assign A_rho[1][3][13]    = A[1][3][32];
    assign A_rho[1][3][14]    = A[1][3][33];
    assign A_rho[1][3][15]    = A[1][3][34];
    assign A_rho[1][3][16]    = A[1][3][35];
    assign A_rho[1][3][17]    = A[1][3][36];
    assign A_rho[1][3][18]    = A[1][3][37];
    assign A_rho[1][3][19]    = A[1][3][38];
    assign A_rho[1][3][20]    = A[1][3][39];
    assign A_rho[1][3][21]    = A[1][3][40];
    assign A_rho[1][3][22]    = A[1][3][41];
    assign A_rho[1][3][23]    = A[1][3][42];
    assign A_rho[1][3][24]    = A[1][3][43];
    assign A_rho[1][3][25]    = A[1][3][44];
    assign A_rho[1][3][26]    = A[1][3][45];
    assign A_rho[1][3][27]    = A[1][3][46];
    assign A_rho[1][3][28]    = A[1][3][47];
    assign A_rho[1][3][29]    = A[1][3][48];
    assign A_rho[1][3][30]    = A[1][3][49];
    assign A_rho[1][3][31]    = A[1][3][50];
    assign A_rho[1][3][32]    = A[1][3][51];
    assign A_rho[1][3][33]    = A[1][3][52];
    assign A_rho[1][3][34]    = A[1][3][53];
    assign A_rho[1][3][35]    = A[1][3][54];
    assign A_rho[1][3][36]    = A[1][3][55];
    assign A_rho[1][3][37]    = A[1][3][56];
    assign A_rho[1][3][38]    = A[1][3][57];
    assign A_rho[1][3][39]    = A[1][3][58];
    assign A_rho[1][3][40]    = A[1][3][59];
    assign A_rho[1][3][41]    = A[1][3][60];
    assign A_rho[1][3][42]    = A[1][3][61];
    assign A_rho[1][3][43]    = A[1][3][62];
    assign A_rho[1][3][44]    = A[1][3][63];
    assign A_rho[1][3][45]    = A[1][3][0];
    assign A_rho[1][3][46]    = A[1][3][1];
    assign A_rho[1][3][47]    = A[1][3][2];
    assign A_rho[1][3][48]    = A[1][3][3];
    assign A_rho[1][3][49]    = A[1][3][4];
    assign A_rho[1][3][50]    = A[1][3][5];
    assign A_rho[1][3][51]    = A[1][3][6];
    assign A_rho[1][3][52]    = A[1][3][7];
    assign A_rho[1][3][53]    = A[1][3][8];
    assign A_rho[1][3][54]    = A[1][3][9];
    assign A_rho[1][3][55]    = A[1][3][10];
    assign A_rho[1][3][56]    = A[1][3][11];
    assign A_rho[1][3][57]    = A[1][3][12];
    assign A_rho[1][3][58]    = A[1][3][13];
    assign A_rho[1][3][59]    = A[1][3][14];
    assign A_rho[1][3][60]    = A[1][3][15];
    assign A_rho[1][3][61]    = A[1][3][16];
    assign A_rho[1][3][62]    = A[1][3][17];
    assign A_rho[1][3][63]    = A[1][3][18];
    assign A_rho[3][1][0]    = A[3][1][9];
    assign A_rho[3][1][1]    = A[3][1][10];
    assign A_rho[3][1][2]    = A[3][1][11];
    assign A_rho[3][1][3]    = A[3][1][12];
    assign A_rho[3][1][4]    = A[3][1][13];
    assign A_rho[3][1][5]    = A[3][1][14];
    assign A_rho[3][1][6]    = A[3][1][15];
    assign A_rho[3][1][7]    = A[3][1][16];
    assign A_rho[3][1][8]    = A[3][1][17];
    assign A_rho[3][1][9]    = A[3][1][18];
    assign A_rho[3][1][10]    = A[3][1][19];
    assign A_rho[3][1][11]    = A[3][1][20];
    assign A_rho[3][1][12]    = A[3][1][21];
    assign A_rho[3][1][13]    = A[3][1][22];
    assign A_rho[3][1][14]    = A[3][1][23];
    assign A_rho[3][1][15]    = A[3][1][24];
    assign A_rho[3][1][16]    = A[3][1][25];
    assign A_rho[3][1][17]    = A[3][1][26];
    assign A_rho[3][1][18]    = A[3][1][27];
    assign A_rho[3][1][19]    = A[3][1][28];
    assign A_rho[3][1][20]    = A[3][1][29];
    assign A_rho[3][1][21]    = A[3][1][30];
    assign A_rho[3][1][22]    = A[3][1][31];
    assign A_rho[3][1][23]    = A[3][1][32];
    assign A_rho[3][1][24]    = A[3][1][33];
    assign A_rho[3][1][25]    = A[3][1][34];
    assign A_rho[3][1][26]    = A[3][1][35];
    assign A_rho[3][1][27]    = A[3][1][36];
    assign A_rho[3][1][28]    = A[3][1][37];
    assign A_rho[3][1][29]    = A[3][1][38];
    assign A_rho[3][1][30]    = A[3][1][39];
    assign A_rho[3][1][31]    = A[3][1][40];
    assign A_rho[3][1][32]    = A[3][1][41];
    assign A_rho[3][1][33]    = A[3][1][42];
    assign A_rho[3][1][34]    = A[3][1][43];
    assign A_rho[3][1][35]    = A[3][1][44];
    assign A_rho[3][1][36]    = A[3][1][45];
    assign A_rho[3][1][37]    = A[3][1][46];
    assign A_rho[3][1][38]    = A[3][1][47];
    assign A_rho[3][1][39]    = A[3][1][48];
    assign A_rho[3][1][40]    = A[3][1][49];
    assign A_rho[3][1][41]    = A[3][1][50];
    assign A_rho[3][1][42]    = A[3][1][51];
    assign A_rho[3][1][43]    = A[3][1][52];
    assign A_rho[3][1][44]    = A[3][1][53];
    assign A_rho[3][1][45]    = A[3][1][54];
    assign A_rho[3][1][46]    = A[3][1][55];
    assign A_rho[3][1][47]    = A[3][1][56];
    assign A_rho[3][1][48]    = A[3][1][57];
    assign A_rho[3][1][49]    = A[3][1][58];
    assign A_rho[3][1][50]    = A[3][1][59];
    assign A_rho[3][1][51]    = A[3][1][60];
    assign A_rho[3][1][52]    = A[3][1][61];
    assign A_rho[3][1][53]    = A[3][1][62];
    assign A_rho[3][1][54]    = A[3][1][63];
    assign A_rho[3][1][55]    = A[3][1][0];
    assign A_rho[3][1][56]    = A[3][1][1];
    assign A_rho[3][1][57]    = A[3][1][2];
    assign A_rho[3][1][58]    = A[3][1][3];
    assign A_rho[3][1][59]    = A[3][1][4];
    assign A_rho[3][1][60]    = A[3][1][5];
    assign A_rho[3][1][61]    = A[3][1][6];
    assign A_rho[3][1][62]    = A[3][1][7];
    assign A_rho[3][1][63]    = A[3][1][8];
    assign A_rho[1][4][0]    = A[1][4][62];
    assign A_rho[1][4][1]    = A[1][4][63];
    assign A_rho[1][4][2]    = A[1][4][0];
    assign A_rho[1][4][3]    = A[1][4][1];
    assign A_rho[1][4][4]    = A[1][4][2];
    assign A_rho[1][4][5]    = A[1][4][3];
    assign A_rho[1][4][6]    = A[1][4][4];
    assign A_rho[1][4][7]    = A[1][4][5];
    assign A_rho[1][4][8]    = A[1][4][6];
    assign A_rho[1][4][9]    = A[1][4][7];
    assign A_rho[1][4][10]    = A[1][4][8];
    assign A_rho[1][4][11]    = A[1][4][9];
    assign A_rho[1][4][12]    = A[1][4][10];
    assign A_rho[1][4][13]    = A[1][4][11];
    assign A_rho[1][4][14]    = A[1][4][12];
    assign A_rho[1][4][15]    = A[1][4][13];
    assign A_rho[1][4][16]    = A[1][4][14];
    assign A_rho[1][4][17]    = A[1][4][15];
    assign A_rho[1][4][18]    = A[1][4][16];
    assign A_rho[1][4][19]    = A[1][4][17];
    assign A_rho[1][4][20]    = A[1][4][18];
    assign A_rho[1][4][21]    = A[1][4][19];
    assign A_rho[1][4][22]    = A[1][4][20];
    assign A_rho[1][4][23]    = A[1][4][21];
    assign A_rho[1][4][24]    = A[1][4][22];
    assign A_rho[1][4][25]    = A[1][4][23];
    assign A_rho[1][4][26]    = A[1][4][24];
    assign A_rho[1][4][27]    = A[1][4][25];
    assign A_rho[1][4][28]    = A[1][4][26];
    assign A_rho[1][4][29]    = A[1][4][27];
    assign A_rho[1][4][30]    = A[1][4][28];
    assign A_rho[1][4][31]    = A[1][4][29];
    assign A_rho[1][4][32]    = A[1][4][30];
    assign A_rho[1][4][33]    = A[1][4][31];
    assign A_rho[1][4][34]    = A[1][4][32];
    assign A_rho[1][4][35]    = A[1][4][33];
    assign A_rho[1][4][36]    = A[1][4][34];
    assign A_rho[1][4][37]    = A[1][4][35];
    assign A_rho[1][4][38]    = A[1][4][36];
    assign A_rho[1][4][39]    = A[1][4][37];
    assign A_rho[1][4][40]    = A[1][4][38];
    assign A_rho[1][4][41]    = A[1][4][39];
    assign A_rho[1][4][42]    = A[1][4][40];
    assign A_rho[1][4][43]    = A[1][4][41];
    assign A_rho[1][4][44]    = A[1][4][42];
    assign A_rho[1][4][45]    = A[1][4][43];
    assign A_rho[1][4][46]    = A[1][4][44];
    assign A_rho[1][4][47]    = A[1][4][45];
    assign A_rho[1][4][48]    = A[1][4][46];
    assign A_rho[1][4][49]    = A[1][4][47];
    assign A_rho[1][4][50]    = A[1][4][48];
    assign A_rho[1][4][51]    = A[1][4][49];
    assign A_rho[1][4][52]    = A[1][4][50];
    assign A_rho[1][4][53]    = A[1][4][51];
    assign A_rho[1][4][54]    = A[1][4][52];
    assign A_rho[1][4][55]    = A[1][4][53];
    assign A_rho[1][4][56]    = A[1][4][54];
    assign A_rho[1][4][57]    = A[1][4][55];
    assign A_rho[1][4][58]    = A[1][4][56];
    assign A_rho[1][4][59]    = A[1][4][57];
    assign A_rho[1][4][60]    = A[1][4][58];
    assign A_rho[1][4][61]    = A[1][4][59];
    assign A_rho[1][4][62]    = A[1][4][60];
    assign A_rho[1][4][63]    = A[1][4][61];
    assign A_rho[4][4][0]    = A[4][4][50];
    assign A_rho[4][4][1]    = A[4][4][51];
    assign A_rho[4][4][2]    = A[4][4][52];
    assign A_rho[4][4][3]    = A[4][4][53];
    assign A_rho[4][4][4]    = A[4][4][54];
    assign A_rho[4][4][5]    = A[4][4][55];
    assign A_rho[4][4][6]    = A[4][4][56];
    assign A_rho[4][4][7]    = A[4][4][57];
    assign A_rho[4][4][8]    = A[4][4][58];
    assign A_rho[4][4][9]    = A[4][4][59];
    assign A_rho[4][4][10]    = A[4][4][60];
    assign A_rho[4][4][11]    = A[4][4][61];
    assign A_rho[4][4][12]    = A[4][4][62];
    assign A_rho[4][4][13]    = A[4][4][63];
    assign A_rho[4][4][14]    = A[4][4][0];
    assign A_rho[4][4][15]    = A[4][4][1];
    assign A_rho[4][4][16]    = A[4][4][2];
    assign A_rho[4][4][17]    = A[4][4][3];
    assign A_rho[4][4][18]    = A[4][4][4];
    assign A_rho[4][4][19]    = A[4][4][5];
    assign A_rho[4][4][20]    = A[4][4][6];
    assign A_rho[4][4][21]    = A[4][4][7];
    assign A_rho[4][4][22]    = A[4][4][8];
    assign A_rho[4][4][23]    = A[4][4][9];
    assign A_rho[4][4][24]    = A[4][4][10];
    assign A_rho[4][4][25]    = A[4][4][11];
    assign A_rho[4][4][26]    = A[4][4][12];
    assign A_rho[4][4][27]    = A[4][4][13];
    assign A_rho[4][4][28]    = A[4][4][14];
    assign A_rho[4][4][29]    = A[4][4][15];
    assign A_rho[4][4][30]    = A[4][4][16];
    assign A_rho[4][4][31]    = A[4][4][17];
    assign A_rho[4][4][32]    = A[4][4][18];
    assign A_rho[4][4][33]    = A[4][4][19];
    assign A_rho[4][4][34]    = A[4][4][20];
    assign A_rho[4][4][35]    = A[4][4][21];
    assign A_rho[4][4][36]    = A[4][4][22];
    assign A_rho[4][4][37]    = A[4][4][23];
    assign A_rho[4][4][38]    = A[4][4][24];
    assign A_rho[4][4][39]    = A[4][4][25];
    assign A_rho[4][4][40]    = A[4][4][26];
    assign A_rho[4][4][41]    = A[4][4][27];
    assign A_rho[4][4][42]    = A[4][4][28];
    assign A_rho[4][4][43]    = A[4][4][29];
    assign A_rho[4][4][44]    = A[4][4][30];
    assign A_rho[4][4][45]    = A[4][4][31];
    assign A_rho[4][4][46]    = A[4][4][32];
    assign A_rho[4][4][47]    = A[4][4][33];
    assign A_rho[4][4][48]    = A[4][4][34];
    assign A_rho[4][4][49]    = A[4][4][35];
    assign A_rho[4][4][50]    = A[4][4][36];
    assign A_rho[4][4][51]    = A[4][4][37];
    assign A_rho[4][4][52]    = A[4][4][38];
    assign A_rho[4][4][53]    = A[4][4][39];
    assign A_rho[4][4][54]    = A[4][4][40];
    assign A_rho[4][4][55]    = A[4][4][41];
    assign A_rho[4][4][56]    = A[4][4][42];
    assign A_rho[4][4][57]    = A[4][4][43];
    assign A_rho[4][4][58]    = A[4][4][44];
    assign A_rho[4][4][59]    = A[4][4][45];
    assign A_rho[4][4][60]    = A[4][4][46];
    assign A_rho[4][4][61]    = A[4][4][47];
    assign A_rho[4][4][62]    = A[4][4][48];
    assign A_rho[4][4][63]    = A[4][4][49];
    assign A_rho[4][0][0]    = A[4][0][37];
    assign A_rho[4][0][1]    = A[4][0][38];
    assign A_rho[4][0][2]    = A[4][0][39];
    assign A_rho[4][0][3]    = A[4][0][40];
    assign A_rho[4][0][4]    = A[4][0][41];
    assign A_rho[4][0][5]    = A[4][0][42];
    assign A_rho[4][0][6]    = A[4][0][43];
    assign A_rho[4][0][7]    = A[4][0][44];
    assign A_rho[4][0][8]    = A[4][0][45];
    assign A_rho[4][0][9]    = A[4][0][46];
    assign A_rho[4][0][10]    = A[4][0][47];
    assign A_rho[4][0][11]    = A[4][0][48];
    assign A_rho[4][0][12]    = A[4][0][49];
    assign A_rho[4][0][13]    = A[4][0][50];
    assign A_rho[4][0][14]    = A[4][0][51];
    assign A_rho[4][0][15]    = A[4][0][52];
    assign A_rho[4][0][16]    = A[4][0][53];
    assign A_rho[4][0][17]    = A[4][0][54];
    assign A_rho[4][0][18]    = A[4][0][55];
    assign A_rho[4][0][19]    = A[4][0][56];
    assign A_rho[4][0][20]    = A[4][0][57];
    assign A_rho[4][0][21]    = A[4][0][58];
    assign A_rho[4][0][22]    = A[4][0][59];
    assign A_rho[4][0][23]    = A[4][0][60];
    assign A_rho[4][0][24]    = A[4][0][61];
    assign A_rho[4][0][25]    = A[4][0][62];
    assign A_rho[4][0][26]    = A[4][0][63];
    assign A_rho[4][0][27]    = A[4][0][0];
    assign A_rho[4][0][28]    = A[4][0][1];
    assign A_rho[4][0][29]    = A[4][0][2];
    assign A_rho[4][0][30]    = A[4][0][3];
    assign A_rho[4][0][31]    = A[4][0][4];
    assign A_rho[4][0][32]    = A[4][0][5];
    assign A_rho[4][0][33]    = A[4][0][6];
    assign A_rho[4][0][34]    = A[4][0][7];
    assign A_rho[4][0][35]    = A[4][0][8];
    assign A_rho[4][0][36]    = A[4][0][9];
    assign A_rho[4][0][37]    = A[4][0][10];
    assign A_rho[4][0][38]    = A[4][0][11];
    assign A_rho[4][0][39]    = A[4][0][12];
    assign A_rho[4][0][40]    = A[4][0][13];
    assign A_rho[4][0][41]    = A[4][0][14];
    assign A_rho[4][0][42]    = A[4][0][15];
    assign A_rho[4][0][43]    = A[4][0][16];
    assign A_rho[4][0][44]    = A[4][0][17];
    assign A_rho[4][0][45]    = A[4][0][18];
    assign A_rho[4][0][46]    = A[4][0][19];
    assign A_rho[4][0][47]    = A[4][0][20];
    assign A_rho[4][0][48]    = A[4][0][21];
    assign A_rho[4][0][49]    = A[4][0][22];
    assign A_rho[4][0][50]    = A[4][0][23];
    assign A_rho[4][0][51]    = A[4][0][24];
    assign A_rho[4][0][52]    = A[4][0][25];
    assign A_rho[4][0][53]    = A[4][0][26];
    assign A_rho[4][0][54]    = A[4][0][27];
    assign A_rho[4][0][55]    = A[4][0][28];
    assign A_rho[4][0][56]    = A[4][0][29];
    assign A_rho[4][0][57]    = A[4][0][30];
    assign A_rho[4][0][58]    = A[4][0][31];
    assign A_rho[4][0][59]    = A[4][0][32];
    assign A_rho[4][0][60]    = A[4][0][33];
    assign A_rho[4][0][61]    = A[4][0][34];
    assign A_rho[4][0][62]    = A[4][0][35];
    assign A_rho[4][0][63]    = A[4][0][36];
    assign A_rho[0][3][0]    = A[0][3][23];
    assign A_rho[0][3][1]    = A[0][3][24];
    assign A_rho[0][3][2]    = A[0][3][25];
    assign A_rho[0][3][3]    = A[0][3][26];
    assign A_rho[0][3][4]    = A[0][3][27];
    assign A_rho[0][3][5]    = A[0][3][28];
    assign A_rho[0][3][6]    = A[0][3][29];
    assign A_rho[0][3][7]    = A[0][3][30];
    assign A_rho[0][3][8]    = A[0][3][31];
    assign A_rho[0][3][9]    = A[0][3][32];
    assign A_rho[0][3][10]    = A[0][3][33];
    assign A_rho[0][3][11]    = A[0][3][34];
    assign A_rho[0][3][12]    = A[0][3][35];
    assign A_rho[0][3][13]    = A[0][3][36];
    assign A_rho[0][3][14]    = A[0][3][37];
    assign A_rho[0][3][15]    = A[0][3][38];
    assign A_rho[0][3][16]    = A[0][3][39];
    assign A_rho[0][3][17]    = A[0][3][40];
    assign A_rho[0][3][18]    = A[0][3][41];
    assign A_rho[0][3][19]    = A[0][3][42];
    assign A_rho[0][3][20]    = A[0][3][43];
    assign A_rho[0][3][21]    = A[0][3][44];
    assign A_rho[0][3][22]    = A[0][3][45];
    assign A_rho[0][3][23]    = A[0][3][46];
    assign A_rho[0][3][24]    = A[0][3][47];
    assign A_rho[0][3][25]    = A[0][3][48];
    assign A_rho[0][3][26]    = A[0][3][49];
    assign A_rho[0][3][27]    = A[0][3][50];
    assign A_rho[0][3][28]    = A[0][3][51];
    assign A_rho[0][3][29]    = A[0][3][52];
    assign A_rho[0][3][30]    = A[0][3][53];
    assign A_rho[0][3][31]    = A[0][3][54];
    assign A_rho[0][3][32]    = A[0][3][55];
    assign A_rho[0][3][33]    = A[0][3][56];
    assign A_rho[0][3][34]    = A[0][3][57];
    assign A_rho[0][3][35]    = A[0][3][58];
    assign A_rho[0][3][36]    = A[0][3][59];
    assign A_rho[0][3][37]    = A[0][3][60];
    assign A_rho[0][3][38]    = A[0][3][61];
    assign A_rho[0][3][39]    = A[0][3][62];
    assign A_rho[0][3][40]    = A[0][3][63];
    assign A_rho[0][3][41]    = A[0][3][0];
    assign A_rho[0][3][42]    = A[0][3][1];
    assign A_rho[0][3][43]    = A[0][3][2];
    assign A_rho[0][3][44]    = A[0][3][3];
    assign A_rho[0][3][45]    = A[0][3][4];
    assign A_rho[0][3][46]    = A[0][3][5];
    assign A_rho[0][3][47]    = A[0][3][6];
    assign A_rho[0][3][48]    = A[0][3][7];
    assign A_rho[0][3][49]    = A[0][3][8];
    assign A_rho[0][3][50]    = A[0][3][9];
    assign A_rho[0][3][51]    = A[0][3][10];
    assign A_rho[0][3][52]    = A[0][3][11];
    assign A_rho[0][3][53]    = A[0][3][12];
    assign A_rho[0][3][54]    = A[0][3][13];
    assign A_rho[0][3][55]    = A[0][3][14];
    assign A_rho[0][3][56]    = A[0][3][15];
    assign A_rho[0][3][57]    = A[0][3][16];
    assign A_rho[0][3][58]    = A[0][3][17];
    assign A_rho[0][3][59]    = A[0][3][18];
    assign A_rho[0][3][60]    = A[0][3][19];
    assign A_rho[0][3][61]    = A[0][3][20];
    assign A_rho[0][3][62]    = A[0][3][21];
    assign A_rho[0][3][63]    = A[0][3][22];
    assign A_rho[3][4][0]    = A[3][4][8];
    assign A_rho[3][4][1]    = A[3][4][9];
    assign A_rho[3][4][2]    = A[3][4][10];
    assign A_rho[3][4][3]    = A[3][4][11];
    assign A_rho[3][4][4]    = A[3][4][12];
    assign A_rho[3][4][5]    = A[3][4][13];
    assign A_rho[3][4][6]    = A[3][4][14];
    assign A_rho[3][4][7]    = A[3][4][15];
    assign A_rho[3][4][8]    = A[3][4][16];
    assign A_rho[3][4][9]    = A[3][4][17];
    assign A_rho[3][4][10]    = A[3][4][18];
    assign A_rho[3][4][11]    = A[3][4][19];
    assign A_rho[3][4][12]    = A[3][4][20];
    assign A_rho[3][4][13]    = A[3][4][21];
    assign A_rho[3][4][14]    = A[3][4][22];
    assign A_rho[3][4][15]    = A[3][4][23];
    assign A_rho[3][4][16]    = A[3][4][24];
    assign A_rho[3][4][17]    = A[3][4][25];
    assign A_rho[3][4][18]    = A[3][4][26];
    assign A_rho[3][4][19]    = A[3][4][27];
    assign A_rho[3][4][20]    = A[3][4][28];
    assign A_rho[3][4][21]    = A[3][4][29];
    assign A_rho[3][4][22]    = A[3][4][30];
    assign A_rho[3][4][23]    = A[3][4][31];
    assign A_rho[3][4][24]    = A[3][4][32];
    assign A_rho[3][4][25]    = A[3][4][33];
    assign A_rho[3][4][26]    = A[3][4][34];
    assign A_rho[3][4][27]    = A[3][4][35];
    assign A_rho[3][4][28]    = A[3][4][36];
    assign A_rho[3][4][29]    = A[3][4][37];
    assign A_rho[3][4][30]    = A[3][4][38];
    assign A_rho[3][4][31]    = A[3][4][39];
    assign A_rho[3][4][32]    = A[3][4][40];
    assign A_rho[3][4][33]    = A[3][4][41];
    assign A_rho[3][4][34]    = A[3][4][42];
    assign A_rho[3][4][35]    = A[3][4][43];
    assign A_rho[3][4][36]    = A[3][4][44];
    assign A_rho[3][4][37]    = A[3][4][45];
    assign A_rho[3][4][38]    = A[3][4][46];
    assign A_rho[3][4][39]    = A[3][4][47];
    assign A_rho[3][4][40]    = A[3][4][48];
    assign A_rho[3][4][41]    = A[3][4][49];
    assign A_rho[3][4][42]    = A[3][4][50];
    assign A_rho[3][4][43]    = A[3][4][51];
    assign A_rho[3][4][44]    = A[3][4][52];
    assign A_rho[3][4][45]    = A[3][4][53];
    assign A_rho[3][4][46]    = A[3][4][54];
    assign A_rho[3][4][47]    = A[3][4][55];
    assign A_rho[3][4][48]    = A[3][4][56];
    assign A_rho[3][4][49]    = A[3][4][57];
    assign A_rho[3][4][50]    = A[3][4][58];
    assign A_rho[3][4][51]    = A[3][4][59];
    assign A_rho[3][4][52]    = A[3][4][60];
    assign A_rho[3][4][53]    = A[3][4][61];
    assign A_rho[3][4][54]    = A[3][4][62];
    assign A_rho[3][4][55]    = A[3][4][63];
    assign A_rho[3][4][56]    = A[3][4][0];
    assign A_rho[3][4][57]    = A[3][4][1];
    assign A_rho[3][4][58]    = A[3][4][2];
    assign A_rho[3][4][59]    = A[3][4][3];
    assign A_rho[3][4][60]    = A[3][4][4];
    assign A_rho[3][4][61]    = A[3][4][5];
    assign A_rho[3][4][62]    = A[3][4][6];
    assign A_rho[3][4][63]    = A[3][4][7];
    assign A_rho[4][3][0]    = A[4][3][56];
    assign A_rho[4][3][1]    = A[4][3][57];
    assign A_rho[4][3][2]    = A[4][3][58];
    assign A_rho[4][3][3]    = A[4][3][59];
    assign A_rho[4][3][4]    = A[4][3][60];
    assign A_rho[4][3][5]    = A[4][3][61];
    assign A_rho[4][3][6]    = A[4][3][62];
    assign A_rho[4][3][7]    = A[4][3][63];
    assign A_rho[4][3][8]    = A[4][3][0];
    assign A_rho[4][3][9]    = A[4][3][1];
    assign A_rho[4][3][10]    = A[4][3][2];
    assign A_rho[4][3][11]    = A[4][3][3];
    assign A_rho[4][3][12]    = A[4][3][4];
    assign A_rho[4][3][13]    = A[4][3][5];
    assign A_rho[4][3][14]    = A[4][3][6];
    assign A_rho[4][3][15]    = A[4][3][7];
    assign A_rho[4][3][16]    = A[4][3][8];
    assign A_rho[4][3][17]    = A[4][3][9];
    assign A_rho[4][3][18]    = A[4][3][10];
    assign A_rho[4][3][19]    = A[4][3][11];
    assign A_rho[4][3][20]    = A[4][3][12];
    assign A_rho[4][3][21]    = A[4][3][13];
    assign A_rho[4][3][22]    = A[4][3][14];
    assign A_rho[4][3][23]    = A[4][3][15];
    assign A_rho[4][3][24]    = A[4][3][16];
    assign A_rho[4][3][25]    = A[4][3][17];
    assign A_rho[4][3][26]    = A[4][3][18];
    assign A_rho[4][3][27]    = A[4][3][19];
    assign A_rho[4][3][28]    = A[4][3][20];
    assign A_rho[4][3][29]    = A[4][3][21];
    assign A_rho[4][3][30]    = A[4][3][22];
    assign A_rho[4][3][31]    = A[4][3][23];
    assign A_rho[4][3][32]    = A[4][3][24];
    assign A_rho[4][3][33]    = A[4][3][25];
    assign A_rho[4][3][34]    = A[4][3][26];
    assign A_rho[4][3][35]    = A[4][3][27];
    assign A_rho[4][3][36]    = A[4][3][28];
    assign A_rho[4][3][37]    = A[4][3][29];
    assign A_rho[4][3][38]    = A[4][3][30];
    assign A_rho[4][3][39]    = A[4][3][31];
    assign A_rho[4][3][40]    = A[4][3][32];
    assign A_rho[4][3][41]    = A[4][3][33];
    assign A_rho[4][3][42]    = A[4][3][34];
    assign A_rho[4][3][43]    = A[4][3][35];
    assign A_rho[4][3][44]    = A[4][3][36];
    assign A_rho[4][3][45]    = A[4][3][37];
    assign A_rho[4][3][46]    = A[4][3][38];
    assign A_rho[4][3][47]    = A[4][3][39];
    assign A_rho[4][3][48]    = A[4][3][40];
    assign A_rho[4][3][49]    = A[4][3][41];
    assign A_rho[4][3][50]    = A[4][3][42];
    assign A_rho[4][3][51]    = A[4][3][43];
    assign A_rho[4][3][52]    = A[4][3][44];
    assign A_rho[4][3][53]    = A[4][3][45];
    assign A_rho[4][3][54]    = A[4][3][46];
    assign A_rho[4][3][55]    = A[4][3][47];
    assign A_rho[4][3][56]    = A[4][3][48];
    assign A_rho[4][3][57]    = A[4][3][49];
    assign A_rho[4][3][58]    = A[4][3][50];
    assign A_rho[4][3][59]    = A[4][3][51];
    assign A_rho[4][3][60]    = A[4][3][52];
    assign A_rho[4][3][61]    = A[4][3][53];
    assign A_rho[4][3][62]    = A[4][3][54];
    assign A_rho[4][3][63]    = A[4][3][55];
    assign A_rho[3][2][0]    = A[3][2][39];
    assign A_rho[3][2][1]    = A[3][2][40];
    assign A_rho[3][2][2]    = A[3][2][41];
    assign A_rho[3][2][3]    = A[3][2][42];
    assign A_rho[3][2][4]    = A[3][2][43];
    assign A_rho[3][2][5]    = A[3][2][44];
    assign A_rho[3][2][6]    = A[3][2][45];
    assign A_rho[3][2][7]    = A[3][2][46];
    assign A_rho[3][2][8]    = A[3][2][47];
    assign A_rho[3][2][9]    = A[3][2][48];
    assign A_rho[3][2][10]    = A[3][2][49];
    assign A_rho[3][2][11]    = A[3][2][50];
    assign A_rho[3][2][12]    = A[3][2][51];
    assign A_rho[3][2][13]    = A[3][2][52];
    assign A_rho[3][2][14]    = A[3][2][53];
    assign A_rho[3][2][15]    = A[3][2][54];
    assign A_rho[3][2][16]    = A[3][2][55];
    assign A_rho[3][2][17]    = A[3][2][56];
    assign A_rho[3][2][18]    = A[3][2][57];
    assign A_rho[3][2][19]    = A[3][2][58];
    assign A_rho[3][2][20]    = A[3][2][59];
    assign A_rho[3][2][21]    = A[3][2][60];
    assign A_rho[3][2][22]    = A[3][2][61];
    assign A_rho[3][2][23]    = A[3][2][62];
    assign A_rho[3][2][24]    = A[3][2][63];
    assign A_rho[3][2][25]    = A[3][2][0];
    assign A_rho[3][2][26]    = A[3][2][1];
    assign A_rho[3][2][27]    = A[3][2][2];
    assign A_rho[3][2][28]    = A[3][2][3];
    assign A_rho[3][2][29]    = A[3][2][4];
    assign A_rho[3][2][30]    = A[3][2][5];
    assign A_rho[3][2][31]    = A[3][2][6];
    assign A_rho[3][2][32]    = A[3][2][7];
    assign A_rho[3][2][33]    = A[3][2][8];
    assign A_rho[3][2][34]    = A[3][2][9];
    assign A_rho[3][2][35]    = A[3][2][10];
    assign A_rho[3][2][36]    = A[3][2][11];
    assign A_rho[3][2][37]    = A[3][2][12];
    assign A_rho[3][2][38]    = A[3][2][13];
    assign A_rho[3][2][39]    = A[3][2][14];
    assign A_rho[3][2][40]    = A[3][2][15];
    assign A_rho[3][2][41]    = A[3][2][16];
    assign A_rho[3][2][42]    = A[3][2][17];
    assign A_rho[3][2][43]    = A[3][2][18];
    assign A_rho[3][2][44]    = A[3][2][19];
    assign A_rho[3][2][45]    = A[3][2][20];
    assign A_rho[3][2][46]    = A[3][2][21];
    assign A_rho[3][2][47]    = A[3][2][22];
    assign A_rho[3][2][48]    = A[3][2][23];
    assign A_rho[3][2][49]    = A[3][2][24];
    assign A_rho[3][2][50]    = A[3][2][25];
    assign A_rho[3][2][51]    = A[3][2][26];
    assign A_rho[3][2][52]    = A[3][2][27];
    assign A_rho[3][2][53]    = A[3][2][28];
    assign A_rho[3][2][54]    = A[3][2][29];
    assign A_rho[3][2][55]    = A[3][2][30];
    assign A_rho[3][2][56]    = A[3][2][31];
    assign A_rho[3][2][57]    = A[3][2][32];
    assign A_rho[3][2][58]    = A[3][2][33];
    assign A_rho[3][2][59]    = A[3][2][34];
    assign A_rho[3][2][60]    = A[3][2][35];
    assign A_rho[3][2][61]    = A[3][2][36];
    assign A_rho[3][2][62]    = A[3][2][37];
    assign A_rho[3][2][63]    = A[3][2][38];
    assign A_rho[2][2][0]    = A[2][2][21];
    assign A_rho[2][2][1]    = A[2][2][22];
    assign A_rho[2][2][2]    = A[2][2][23];
    assign A_rho[2][2][3]    = A[2][2][24];
    assign A_rho[2][2][4]    = A[2][2][25];
    assign A_rho[2][2][5]    = A[2][2][26];
    assign A_rho[2][2][6]    = A[2][2][27];
    assign A_rho[2][2][7]    = A[2][2][28];
    assign A_rho[2][2][8]    = A[2][2][29];
    assign A_rho[2][2][9]    = A[2][2][30];
    assign A_rho[2][2][10]    = A[2][2][31];
    assign A_rho[2][2][11]    = A[2][2][32];
    assign A_rho[2][2][12]    = A[2][2][33];
    assign A_rho[2][2][13]    = A[2][2][34];
    assign A_rho[2][2][14]    = A[2][2][35];
    assign A_rho[2][2][15]    = A[2][2][36];
    assign A_rho[2][2][16]    = A[2][2][37];
    assign A_rho[2][2][17]    = A[2][2][38];
    assign A_rho[2][2][18]    = A[2][2][39];
    assign A_rho[2][2][19]    = A[2][2][40];
    assign A_rho[2][2][20]    = A[2][2][41];
    assign A_rho[2][2][21]    = A[2][2][42];
    assign A_rho[2][2][22]    = A[2][2][43];
    assign A_rho[2][2][23]    = A[2][2][44];
    assign A_rho[2][2][24]    = A[2][2][45];
    assign A_rho[2][2][25]    = A[2][2][46];
    assign A_rho[2][2][26]    = A[2][2][47];
    assign A_rho[2][2][27]    = A[2][2][48];
    assign A_rho[2][2][28]    = A[2][2][49];
    assign A_rho[2][2][29]    = A[2][2][50];
    assign A_rho[2][2][30]    = A[2][2][51];
    assign A_rho[2][2][31]    = A[2][2][52];
    assign A_rho[2][2][32]    = A[2][2][53];
    assign A_rho[2][2][33]    = A[2][2][54];
    assign A_rho[2][2][34]    = A[2][2][55];
    assign A_rho[2][2][35]    = A[2][2][56];
    assign A_rho[2][2][36]    = A[2][2][57];
    assign A_rho[2][2][37]    = A[2][2][58];
    assign A_rho[2][2][38]    = A[2][2][59];
    assign A_rho[2][2][39]    = A[2][2][60];
    assign A_rho[2][2][40]    = A[2][2][61];
    assign A_rho[2][2][41]    = A[2][2][62];
    assign A_rho[2][2][42]    = A[2][2][63];
    assign A_rho[2][2][43]    = A[2][2][0];
    assign A_rho[2][2][44]    = A[2][2][1];
    assign A_rho[2][2][45]    = A[2][2][2];
    assign A_rho[2][2][46]    = A[2][2][3];
    assign A_rho[2][2][47]    = A[2][2][4];
    assign A_rho[2][2][48]    = A[2][2][5];
    assign A_rho[2][2][49]    = A[2][2][6];
    assign A_rho[2][2][50]    = A[2][2][7];
    assign A_rho[2][2][51]    = A[2][2][8];
    assign A_rho[2][2][52]    = A[2][2][9];
    assign A_rho[2][2][53]    = A[2][2][10];
    assign A_rho[2][2][54]    = A[2][2][11];
    assign A_rho[2][2][55]    = A[2][2][12];
    assign A_rho[2][2][56]    = A[2][2][13];
    assign A_rho[2][2][57]    = A[2][2][14];
    assign A_rho[2][2][58]    = A[2][2][15];
    assign A_rho[2][2][59]    = A[2][2][16];
    assign A_rho[2][2][60]    = A[2][2][17];
    assign A_rho[2][2][61]    = A[2][2][18];
    assign A_rho[2][2][62]    = A[2][2][19];
    assign A_rho[2][2][63]    = A[2][2][20];
    assign A_rho[2][0][0]    = A[2][0][2];
    assign A_rho[2][0][1]    = A[2][0][3];
    assign A_rho[2][0][2]    = A[2][0][4];
    assign A_rho[2][0][3]    = A[2][0][5];
    assign A_rho[2][0][4]    = A[2][0][6];
    assign A_rho[2][0][5]    = A[2][0][7];
    assign A_rho[2][0][6]    = A[2][0][8];
    assign A_rho[2][0][7]    = A[2][0][9];
    assign A_rho[2][0][8]    = A[2][0][10];
    assign A_rho[2][0][9]    = A[2][0][11];
    assign A_rho[2][0][10]    = A[2][0][12];
    assign A_rho[2][0][11]    = A[2][0][13];
    assign A_rho[2][0][12]    = A[2][0][14];
    assign A_rho[2][0][13]    = A[2][0][15];
    assign A_rho[2][0][14]    = A[2][0][16];
    assign A_rho[2][0][15]    = A[2][0][17];
    assign A_rho[2][0][16]    = A[2][0][18];
    assign A_rho[2][0][17]    = A[2][0][19];
    assign A_rho[2][0][18]    = A[2][0][20];
    assign A_rho[2][0][19]    = A[2][0][21];
    assign A_rho[2][0][20]    = A[2][0][22];
    assign A_rho[2][0][21]    = A[2][0][23];
    assign A_rho[2][0][22]    = A[2][0][24];
    assign A_rho[2][0][23]    = A[2][0][25];
    assign A_rho[2][0][24]    = A[2][0][26];
    assign A_rho[2][0][25]    = A[2][0][27];
    assign A_rho[2][0][26]    = A[2][0][28];
    assign A_rho[2][0][27]    = A[2][0][29];
    assign A_rho[2][0][28]    = A[2][0][30];
    assign A_rho[2][0][29]    = A[2][0][31];
    assign A_rho[2][0][30]    = A[2][0][32];
    assign A_rho[2][0][31]    = A[2][0][33];
    assign A_rho[2][0][32]    = A[2][0][34];
    assign A_rho[2][0][33]    = A[2][0][35];
    assign A_rho[2][0][34]    = A[2][0][36];
    assign A_rho[2][0][35]    = A[2][0][37];
    assign A_rho[2][0][36]    = A[2][0][38];
    assign A_rho[2][0][37]    = A[2][0][39];
    assign A_rho[2][0][38]    = A[2][0][40];
    assign A_rho[2][0][39]    = A[2][0][41];
    assign A_rho[2][0][40]    = A[2][0][42];
    assign A_rho[2][0][41]    = A[2][0][43];
    assign A_rho[2][0][42]    = A[2][0][44];
    assign A_rho[2][0][43]    = A[2][0][45];
    assign A_rho[2][0][44]    = A[2][0][46];
    assign A_rho[2][0][45]    = A[2][0][47];
    assign A_rho[2][0][46]    = A[2][0][48];
    assign A_rho[2][0][47]    = A[2][0][49];
    assign A_rho[2][0][48]    = A[2][0][50];
    assign A_rho[2][0][49]    = A[2][0][51];
    assign A_rho[2][0][50]    = A[2][0][52];
    assign A_rho[2][0][51]    = A[2][0][53];
    assign A_rho[2][0][52]    = A[2][0][54];
    assign A_rho[2][0][53]    = A[2][0][55];
    assign A_rho[2][0][54]    = A[2][0][56];
    assign A_rho[2][0][55]    = A[2][0][57];
    assign A_rho[2][0][56]    = A[2][0][58];
    assign A_rho[2][0][57]    = A[2][0][59];
    assign A_rho[2][0][58]    = A[2][0][60];
    assign A_rho[2][0][59]    = A[2][0][61];
    assign A_rho[2][0][60]    = A[2][0][62];
    assign A_rho[2][0][61]    = A[2][0][63];
    assign A_rho[2][0][62]    = A[2][0][0];
    assign A_rho[2][0][63]    = A[2][0][1];
    assign A_rho[0][4][0]    = A[0][4][46];
    assign A_rho[0][4][1]    = A[0][4][47];
    assign A_rho[0][4][2]    = A[0][4][48];
    assign A_rho[0][4][3]    = A[0][4][49];
    assign A_rho[0][4][4]    = A[0][4][50];
    assign A_rho[0][4][5]    = A[0][4][51];
    assign A_rho[0][4][6]    = A[0][4][52];
    assign A_rho[0][4][7]    = A[0][4][53];
    assign A_rho[0][4][8]    = A[0][4][54];
    assign A_rho[0][4][9]    = A[0][4][55];
    assign A_rho[0][4][10]    = A[0][4][56];
    assign A_rho[0][4][11]    = A[0][4][57];
    assign A_rho[0][4][12]    = A[0][4][58];
    assign A_rho[0][4][13]    = A[0][4][59];
    assign A_rho[0][4][14]    = A[0][4][60];
    assign A_rho[0][4][15]    = A[0][4][61];
    assign A_rho[0][4][16]    = A[0][4][62];
    assign A_rho[0][4][17]    = A[0][4][63];
    assign A_rho[0][4][18]    = A[0][4][0];
    assign A_rho[0][4][19]    = A[0][4][1];
    assign A_rho[0][4][20]    = A[0][4][2];
    assign A_rho[0][4][21]    = A[0][4][3];
    assign A_rho[0][4][22]    = A[0][4][4];
    assign A_rho[0][4][23]    = A[0][4][5];
    assign A_rho[0][4][24]    = A[0][4][6];
    assign A_rho[0][4][25]    = A[0][4][7];
    assign A_rho[0][4][26]    = A[0][4][8];
    assign A_rho[0][4][27]    = A[0][4][9];
    assign A_rho[0][4][28]    = A[0][4][10];
    assign A_rho[0][4][29]    = A[0][4][11];
    assign A_rho[0][4][30]    = A[0][4][12];
    assign A_rho[0][4][31]    = A[0][4][13];
    assign A_rho[0][4][32]    = A[0][4][14];
    assign A_rho[0][4][33]    = A[0][4][15];
    assign A_rho[0][4][34]    = A[0][4][16];
    assign A_rho[0][4][35]    = A[0][4][17];
    assign A_rho[0][4][36]    = A[0][4][18];
    assign A_rho[0][4][37]    = A[0][4][19];
    assign A_rho[0][4][38]    = A[0][4][20];
    assign A_rho[0][4][39]    = A[0][4][21];
    assign A_rho[0][4][40]    = A[0][4][22];
    assign A_rho[0][4][41]    = A[0][4][23];
    assign A_rho[0][4][42]    = A[0][4][24];
    assign A_rho[0][4][43]    = A[0][4][25];
    assign A_rho[0][4][44]    = A[0][4][26];
    assign A_rho[0][4][45]    = A[0][4][27];
    assign A_rho[0][4][46]    = A[0][4][28];
    assign A_rho[0][4][47]    = A[0][4][29];
    assign A_rho[0][4][48]    = A[0][4][30];
    assign A_rho[0][4][49]    = A[0][4][31];
    assign A_rho[0][4][50]    = A[0][4][32];
    assign A_rho[0][4][51]    = A[0][4][33];
    assign A_rho[0][4][52]    = A[0][4][34];
    assign A_rho[0][4][53]    = A[0][4][35];
    assign A_rho[0][4][54]    = A[0][4][36];
    assign A_rho[0][4][55]    = A[0][4][37];
    assign A_rho[0][4][56]    = A[0][4][38];
    assign A_rho[0][4][57]    = A[0][4][39];
    assign A_rho[0][4][58]    = A[0][4][40];
    assign A_rho[0][4][59]    = A[0][4][41];
    assign A_rho[0][4][60]    = A[0][4][42];
    assign A_rho[0][4][61]    = A[0][4][43];
    assign A_rho[0][4][62]    = A[0][4][44];
    assign A_rho[0][4][63]    = A[0][4][45];
    assign A_rho[4][2][0]    = A[4][2][25];
    assign A_rho[4][2][1]    = A[4][2][26];
    assign A_rho[4][2][2]    = A[4][2][27];
    assign A_rho[4][2][3]    = A[4][2][28];
    assign A_rho[4][2][4]    = A[4][2][29];
    assign A_rho[4][2][5]    = A[4][2][30];
    assign A_rho[4][2][6]    = A[4][2][31];
    assign A_rho[4][2][7]    = A[4][2][32];
    assign A_rho[4][2][8]    = A[4][2][33];
    assign A_rho[4][2][9]    = A[4][2][34];
    assign A_rho[4][2][10]    = A[4][2][35];
    assign A_rho[4][2][11]    = A[4][2][36];
    assign A_rho[4][2][12]    = A[4][2][37];
    assign A_rho[4][2][13]    = A[4][2][38];
    assign A_rho[4][2][14]    = A[4][2][39];
    assign A_rho[4][2][15]    = A[4][2][40];
    assign A_rho[4][2][16]    = A[4][2][41];
    assign A_rho[4][2][17]    = A[4][2][42];
    assign A_rho[4][2][18]    = A[4][2][43];
    assign A_rho[4][2][19]    = A[4][2][44];
    assign A_rho[4][2][20]    = A[4][2][45];
    assign A_rho[4][2][21]    = A[4][2][46];
    assign A_rho[4][2][22]    = A[4][2][47];
    assign A_rho[4][2][23]    = A[4][2][48];
    assign A_rho[4][2][24]    = A[4][2][49];
    assign A_rho[4][2][25]    = A[4][2][50];
    assign A_rho[4][2][26]    = A[4][2][51];
    assign A_rho[4][2][27]    = A[4][2][52];
    assign A_rho[4][2][28]    = A[4][2][53];
    assign A_rho[4][2][29]    = A[4][2][54];
    assign A_rho[4][2][30]    = A[4][2][55];
    assign A_rho[4][2][31]    = A[4][2][56];
    assign A_rho[4][2][32]    = A[4][2][57];
    assign A_rho[4][2][33]    = A[4][2][58];
    assign A_rho[4][2][34]    = A[4][2][59];
    assign A_rho[4][2][35]    = A[4][2][60];
    assign A_rho[4][2][36]    = A[4][2][61];
    assign A_rho[4][2][37]    = A[4][2][62];
    assign A_rho[4][2][38]    = A[4][2][63];
    assign A_rho[4][2][39]    = A[4][2][0];
    assign A_rho[4][2][40]    = A[4][2][1];
    assign A_rho[4][2][41]    = A[4][2][2];
    assign A_rho[4][2][42]    = A[4][2][3];
    assign A_rho[4][2][43]    = A[4][2][4];
    assign A_rho[4][2][44]    = A[4][2][5];
    assign A_rho[4][2][45]    = A[4][2][6];
    assign A_rho[4][2][46]    = A[4][2][7];
    assign A_rho[4][2][47]    = A[4][2][8];
    assign A_rho[4][2][48]    = A[4][2][9];
    assign A_rho[4][2][49]    = A[4][2][10];
    assign A_rho[4][2][50]    = A[4][2][11];
    assign A_rho[4][2][51]    = A[4][2][12];
    assign A_rho[4][2][52]    = A[4][2][13];
    assign A_rho[4][2][53]    = A[4][2][14];
    assign A_rho[4][2][54]    = A[4][2][15];
    assign A_rho[4][2][55]    = A[4][2][16];
    assign A_rho[4][2][56]    = A[4][2][17];
    assign A_rho[4][2][57]    = A[4][2][18];
    assign A_rho[4][2][58]    = A[4][2][19];
    assign A_rho[4][2][59]    = A[4][2][20];
    assign A_rho[4][2][60]    = A[4][2][21];
    assign A_rho[4][2][61]    = A[4][2][22];
    assign A_rho[4][2][62]    = A[4][2][23];
    assign A_rho[4][2][63]    = A[4][2][24];
    assign A_rho[2][4][0]    = A[2][4][3];
    assign A_rho[2][4][1]    = A[2][4][4];
    assign A_rho[2][4][2]    = A[2][4][5];
    assign A_rho[2][4][3]    = A[2][4][6];
    assign A_rho[2][4][4]    = A[2][4][7];
    assign A_rho[2][4][5]    = A[2][4][8];
    assign A_rho[2][4][6]    = A[2][4][9];
    assign A_rho[2][4][7]    = A[2][4][10];
    assign A_rho[2][4][8]    = A[2][4][11];
    assign A_rho[2][4][9]    = A[2][4][12];
    assign A_rho[2][4][10]    = A[2][4][13];
    assign A_rho[2][4][11]    = A[2][4][14];
    assign A_rho[2][4][12]    = A[2][4][15];
    assign A_rho[2][4][13]    = A[2][4][16];
    assign A_rho[2][4][14]    = A[2][4][17];
    assign A_rho[2][4][15]    = A[2][4][18];
    assign A_rho[2][4][16]    = A[2][4][19];
    assign A_rho[2][4][17]    = A[2][4][20];
    assign A_rho[2][4][18]    = A[2][4][21];
    assign A_rho[2][4][19]    = A[2][4][22];
    assign A_rho[2][4][20]    = A[2][4][23];
    assign A_rho[2][4][21]    = A[2][4][24];
    assign A_rho[2][4][22]    = A[2][4][25];
    assign A_rho[2][4][23]    = A[2][4][26];
    assign A_rho[2][4][24]    = A[2][4][27];
    assign A_rho[2][4][25]    = A[2][4][28];
    assign A_rho[2][4][26]    = A[2][4][29];
    assign A_rho[2][4][27]    = A[2][4][30];
    assign A_rho[2][4][28]    = A[2][4][31];
    assign A_rho[2][4][29]    = A[2][4][32];
    assign A_rho[2][4][30]    = A[2][4][33];
    assign A_rho[2][4][31]    = A[2][4][34];
    assign A_rho[2][4][32]    = A[2][4][35];
    assign A_rho[2][4][33]    = A[2][4][36];
    assign A_rho[2][4][34]    = A[2][4][37];
    assign A_rho[2][4][35]    = A[2][4][38];
    assign A_rho[2][4][36]    = A[2][4][39];
    assign A_rho[2][4][37]    = A[2][4][40];
    assign A_rho[2][4][38]    = A[2][4][41];
    assign A_rho[2][4][39]    = A[2][4][42];
    assign A_rho[2][4][40]    = A[2][4][43];
    assign A_rho[2][4][41]    = A[2][4][44];
    assign A_rho[2][4][42]    = A[2][4][45];
    assign A_rho[2][4][43]    = A[2][4][46];
    assign A_rho[2][4][44]    = A[2][4][47];
    assign A_rho[2][4][45]    = A[2][4][48];
    assign A_rho[2][4][46]    = A[2][4][49];
    assign A_rho[2][4][47]    = A[2][4][50];
    assign A_rho[2][4][48]    = A[2][4][51];
    assign A_rho[2][4][49]    = A[2][4][52];
    assign A_rho[2][4][50]    = A[2][4][53];
    assign A_rho[2][4][51]    = A[2][4][54];
    assign A_rho[2][4][52]    = A[2][4][55];
    assign A_rho[2][4][53]    = A[2][4][56];
    assign A_rho[2][4][54]    = A[2][4][57];
    assign A_rho[2][4][55]    = A[2][4][58];
    assign A_rho[2][4][56]    = A[2][4][59];
    assign A_rho[2][4][57]    = A[2][4][60];
    assign A_rho[2][4][58]    = A[2][4][61];
    assign A_rho[2][4][59]    = A[2][4][62];
    assign A_rho[2][4][60]    = A[2][4][63];
    assign A_rho[2][4][61]    = A[2][4][0];
    assign A_rho[2][4][62]    = A[2][4][1];
    assign A_rho[2][4][63]    = A[2][4][2];
    assign A_rho[4][1][0]    = A[4][1][44];
    assign A_rho[4][1][1]    = A[4][1][45];
    assign A_rho[4][1][2]    = A[4][1][46];
    assign A_rho[4][1][3]    = A[4][1][47];
    assign A_rho[4][1][4]    = A[4][1][48];
    assign A_rho[4][1][5]    = A[4][1][49];
    assign A_rho[4][1][6]    = A[4][1][50];
    assign A_rho[4][1][7]    = A[4][1][51];
    assign A_rho[4][1][8]    = A[4][1][52];
    assign A_rho[4][1][9]    = A[4][1][53];
    assign A_rho[4][1][10]    = A[4][1][54];
    assign A_rho[4][1][11]    = A[4][1][55];
    assign A_rho[4][1][12]    = A[4][1][56];
    assign A_rho[4][1][13]    = A[4][1][57];
    assign A_rho[4][1][14]    = A[4][1][58];
    assign A_rho[4][1][15]    = A[4][1][59];
    assign A_rho[4][1][16]    = A[4][1][60];
    assign A_rho[4][1][17]    = A[4][1][61];
    assign A_rho[4][1][18]    = A[4][1][62];
    assign A_rho[4][1][19]    = A[4][1][63];
    assign A_rho[4][1][20]    = A[4][1][0];
    assign A_rho[4][1][21]    = A[4][1][1];
    assign A_rho[4][1][22]    = A[4][1][2];
    assign A_rho[4][1][23]    = A[4][1][3];
    assign A_rho[4][1][24]    = A[4][1][4];
    assign A_rho[4][1][25]    = A[4][1][5];
    assign A_rho[4][1][26]    = A[4][1][6];
    assign A_rho[4][1][27]    = A[4][1][7];
    assign A_rho[4][1][28]    = A[4][1][8];
    assign A_rho[4][1][29]    = A[4][1][9];
    assign A_rho[4][1][30]    = A[4][1][10];
    assign A_rho[4][1][31]    = A[4][1][11];
    assign A_rho[4][1][32]    = A[4][1][12];
    assign A_rho[4][1][33]    = A[4][1][13];
    assign A_rho[4][1][34]    = A[4][1][14];
    assign A_rho[4][1][35]    = A[4][1][15];
    assign A_rho[4][1][36]    = A[4][1][16];
    assign A_rho[4][1][37]    = A[4][1][17];
    assign A_rho[4][1][38]    = A[4][1][18];
    assign A_rho[4][1][39]    = A[4][1][19];
    assign A_rho[4][1][40]    = A[4][1][20];
    assign A_rho[4][1][41]    = A[4][1][21];
    assign A_rho[4][1][42]    = A[4][1][22];
    assign A_rho[4][1][43]    = A[4][1][23];
    assign A_rho[4][1][44]    = A[4][1][24];
    assign A_rho[4][1][45]    = A[4][1][25];
    assign A_rho[4][1][46]    = A[4][1][26];
    assign A_rho[4][1][47]    = A[4][1][27];
    assign A_rho[4][1][48]    = A[4][1][28];
    assign A_rho[4][1][49]    = A[4][1][29];
    assign A_rho[4][1][50]    = A[4][1][30];
    assign A_rho[4][1][51]    = A[4][1][31];
    assign A_rho[4][1][52]    = A[4][1][32];
    assign A_rho[4][1][53]    = A[4][1][33];
    assign A_rho[4][1][54]    = A[4][1][34];
    assign A_rho[4][1][55]    = A[4][1][35];
    assign A_rho[4][1][56]    = A[4][1][36];
    assign A_rho[4][1][57]    = A[4][1][37];
    assign A_rho[4][1][58]    = A[4][1][38];
    assign A_rho[4][1][59]    = A[4][1][39];
    assign A_rho[4][1][60]    = A[4][1][40];
    assign A_rho[4][1][61]    = A[4][1][41];
    assign A_rho[4][1][62]    = A[4][1][42];
    assign A_rho[4][1][63]    = A[4][1][43];
    assign A_rho[1][1][0]    = A[1][1][20];
    assign A_rho[1][1][1]    = A[1][1][21];
    assign A_rho[1][1][2]    = A[1][1][22];
    assign A_rho[1][1][3]    = A[1][1][23];
    assign A_rho[1][1][4]    = A[1][1][24];
    assign A_rho[1][1][5]    = A[1][1][25];
    assign A_rho[1][1][6]    = A[1][1][26];
    assign A_rho[1][1][7]    = A[1][1][27];
    assign A_rho[1][1][8]    = A[1][1][28];
    assign A_rho[1][1][9]    = A[1][1][29];
    assign A_rho[1][1][10]    = A[1][1][30];
    assign A_rho[1][1][11]    = A[1][1][31];
    assign A_rho[1][1][12]    = A[1][1][32];
    assign A_rho[1][1][13]    = A[1][1][33];
    assign A_rho[1][1][14]    = A[1][1][34];
    assign A_rho[1][1][15]    = A[1][1][35];
    assign A_rho[1][1][16]    = A[1][1][36];
    assign A_rho[1][1][17]    = A[1][1][37];
    assign A_rho[1][1][18]    = A[1][1][38];
    assign A_rho[1][1][19]    = A[1][1][39];
    assign A_rho[1][1][20]    = A[1][1][40];
    assign A_rho[1][1][21]    = A[1][1][41];
    assign A_rho[1][1][22]    = A[1][1][42];
    assign A_rho[1][1][23]    = A[1][1][43];
    assign A_rho[1][1][24]    = A[1][1][44];
    assign A_rho[1][1][25]    = A[1][1][45];
    assign A_rho[1][1][26]    = A[1][1][46];
    assign A_rho[1][1][27]    = A[1][1][47];
    assign A_rho[1][1][28]    = A[1][1][48];
    assign A_rho[1][1][29]    = A[1][1][49];
    assign A_rho[1][1][30]    = A[1][1][50];
    assign A_rho[1][1][31]    = A[1][1][51];
    assign A_rho[1][1][32]    = A[1][1][52];
    assign A_rho[1][1][33]    = A[1][1][53];
    assign A_rho[1][1][34]    = A[1][1][54];
    assign A_rho[1][1][35]    = A[1][1][55];
    assign A_rho[1][1][36]    = A[1][1][56];
    assign A_rho[1][1][37]    = A[1][1][57];
    assign A_rho[1][1][38]    = A[1][1][58];
    assign A_rho[1][1][39]    = A[1][1][59];
    assign A_rho[1][1][40]    = A[1][1][60];
    assign A_rho[1][1][41]    = A[1][1][61];
    assign A_rho[1][1][42]    = A[1][1][62];
    assign A_rho[1][1][43]    = A[1][1][63];
    assign A_rho[1][1][44]    = A[1][1][0];
    assign A_rho[1][1][45]    = A[1][1][1];
    assign A_rho[1][1][46]    = A[1][1][2];
    assign A_rho[1][1][47]    = A[1][1][3];
    assign A_rho[1][1][48]    = A[1][1][4];
    assign A_rho[1][1][49]    = A[1][1][5];
    assign A_rho[1][1][50]    = A[1][1][6];
    assign A_rho[1][1][51]    = A[1][1][7];
    assign A_rho[1][1][52]    = A[1][1][8];
    assign A_rho[1][1][53]    = A[1][1][9];
    assign A_rho[1][1][54]    = A[1][1][10];
    assign A_rho[1][1][55]    = A[1][1][11];
    assign A_rho[1][1][56]    = A[1][1][12];
    assign A_rho[1][1][57]    = A[1][1][13];
    assign A_rho[1][1][58]    = A[1][1][14];
    assign A_rho[1][1][59]    = A[1][1][15];
    assign A_rho[1][1][60]    = A[1][1][16];
    assign A_rho[1][1][61]    = A[1][1][17];
    assign A_rho[1][1][62]    = A[1][1][18];
    assign A_rho[1][1][63]    = A[1][1][19];
//--------------------------- PI ---------------------------
   assign A_pi[0][0][0]  = A_rho[0][0][0];
   assign A_pi[0][0][1]  = A_rho[0][0][1];
   assign A_pi[0][0][2]  = A_rho[0][0][2];
   assign A_pi[0][0][3]  = A_rho[0][0][3];
   assign A_pi[0][0][4]  = A_rho[0][0][4];
   assign A_pi[0][0][5]  = A_rho[0][0][5];
   assign A_pi[0][0][6]  = A_rho[0][0][6];
   assign A_pi[0][0][7]  = A_rho[0][0][7];
   assign A_pi[0][0][8]  = A_rho[0][0][8];
   assign A_pi[0][0][9]  = A_rho[0][0][9];
   assign A_pi[0][0][10]  = A_rho[0][0][10];
   assign A_pi[0][0][11]  = A_rho[0][0][11];
   assign A_pi[0][0][12]  = A_rho[0][0][12];
   assign A_pi[0][0][13]  = A_rho[0][0][13];
   assign A_pi[0][0][14]  = A_rho[0][0][14];
   assign A_pi[0][0][15]  = A_rho[0][0][15];
   assign A_pi[0][0][16]  = A_rho[0][0][16];
   assign A_pi[0][0][17]  = A_rho[0][0][17];
   assign A_pi[0][0][18]  = A_rho[0][0][18];
   assign A_pi[0][0][19]  = A_rho[0][0][19];
   assign A_pi[0][0][20]  = A_rho[0][0][20];
   assign A_pi[0][0][21]  = A_rho[0][0][21];
   assign A_pi[0][0][22]  = A_rho[0][0][22];
   assign A_pi[0][0][23]  = A_rho[0][0][23];
   assign A_pi[0][0][24]  = A_rho[0][0][24];
   assign A_pi[0][0][25]  = A_rho[0][0][25];
   assign A_pi[0][0][26]  = A_rho[0][0][26];
   assign A_pi[0][0][27]  = A_rho[0][0][27];
   assign A_pi[0][0][28]  = A_rho[0][0][28];
   assign A_pi[0][0][29]  = A_rho[0][0][29];
   assign A_pi[0][0][30]  = A_rho[0][0][30];
   assign A_pi[0][0][31]  = A_rho[0][0][31];
   assign A_pi[0][0][32]  = A_rho[0][0][32];
   assign A_pi[0][0][33]  = A_rho[0][0][33];
   assign A_pi[0][0][34]  = A_rho[0][0][34];
   assign A_pi[0][0][35]  = A_rho[0][0][35];
   assign A_pi[0][0][36]  = A_rho[0][0][36];
   assign A_pi[0][0][37]  = A_rho[0][0][37];
   assign A_pi[0][0][38]  = A_rho[0][0][38];
   assign A_pi[0][0][39]  = A_rho[0][0][39];
   assign A_pi[0][0][40]  = A_rho[0][0][40];
   assign A_pi[0][0][41]  = A_rho[0][0][41];
   assign A_pi[0][0][42]  = A_rho[0][0][42];
   assign A_pi[0][0][43]  = A_rho[0][0][43];
   assign A_pi[0][0][44]  = A_rho[0][0][44];
   assign A_pi[0][0][45]  = A_rho[0][0][45];
   assign A_pi[0][0][46]  = A_rho[0][0][46];
   assign A_pi[0][0][47]  = A_rho[0][0][47];
   assign A_pi[0][0][48]  = A_rho[0][0][48];
   assign A_pi[0][0][49]  = A_rho[0][0][49];
   assign A_pi[0][0][50]  = A_rho[0][0][50];
   assign A_pi[0][0][51]  = A_rho[0][0][51];
   assign A_pi[0][0][52]  = A_rho[0][0][52];
   assign A_pi[0][0][53]  = A_rho[0][0][53];
   assign A_pi[0][0][54]  = A_rho[0][0][54];
   assign A_pi[0][0][55]  = A_rho[0][0][55];
   assign A_pi[0][0][56]  = A_rho[0][0][56];
   assign A_pi[0][0][57]  = A_rho[0][0][57];
   assign A_pi[0][0][58]  = A_rho[0][0][58];
   assign A_pi[0][0][59]  = A_rho[0][0][59];
   assign A_pi[0][0][60]  = A_rho[0][0][60];
   assign A_pi[0][0][61]  = A_rho[0][0][61];
   assign A_pi[0][0][62]  = A_rho[0][0][62];
   assign A_pi[0][0][63]  = A_rho[0][0][63];
   assign A_pi[0][1][0]  = A_rho[3][0][0];
   assign A_pi[0][1][1]  = A_rho[3][0][1];
   assign A_pi[0][1][2]  = A_rho[3][0][2];
   assign A_pi[0][1][3]  = A_rho[3][0][3];
   assign A_pi[0][1][4]  = A_rho[3][0][4];
   assign A_pi[0][1][5]  = A_rho[3][0][5];
   assign A_pi[0][1][6]  = A_rho[3][0][6];
   assign A_pi[0][1][7]  = A_rho[3][0][7];
   assign A_pi[0][1][8]  = A_rho[3][0][8];
   assign A_pi[0][1][9]  = A_rho[3][0][9];
   assign A_pi[0][1][10]  = A_rho[3][0][10];
   assign A_pi[0][1][11]  = A_rho[3][0][11];
   assign A_pi[0][1][12]  = A_rho[3][0][12];
   assign A_pi[0][1][13]  = A_rho[3][0][13];
   assign A_pi[0][1][14]  = A_rho[3][0][14];
   assign A_pi[0][1][15]  = A_rho[3][0][15];
   assign A_pi[0][1][16]  = A_rho[3][0][16];
   assign A_pi[0][1][17]  = A_rho[3][0][17];
   assign A_pi[0][1][18]  = A_rho[3][0][18];
   assign A_pi[0][1][19]  = A_rho[3][0][19];
   assign A_pi[0][1][20]  = A_rho[3][0][20];
   assign A_pi[0][1][21]  = A_rho[3][0][21];
   assign A_pi[0][1][22]  = A_rho[3][0][22];
   assign A_pi[0][1][23]  = A_rho[3][0][23];
   assign A_pi[0][1][24]  = A_rho[3][0][24];
   assign A_pi[0][1][25]  = A_rho[3][0][25];
   assign A_pi[0][1][26]  = A_rho[3][0][26];
   assign A_pi[0][1][27]  = A_rho[3][0][27];
   assign A_pi[0][1][28]  = A_rho[3][0][28];
   assign A_pi[0][1][29]  = A_rho[3][0][29];
   assign A_pi[0][1][30]  = A_rho[3][0][30];
   assign A_pi[0][1][31]  = A_rho[3][0][31];
   assign A_pi[0][1][32]  = A_rho[3][0][32];
   assign A_pi[0][1][33]  = A_rho[3][0][33];
   assign A_pi[0][1][34]  = A_rho[3][0][34];
   assign A_pi[0][1][35]  = A_rho[3][0][35];
   assign A_pi[0][1][36]  = A_rho[3][0][36];
   assign A_pi[0][1][37]  = A_rho[3][0][37];
   assign A_pi[0][1][38]  = A_rho[3][0][38];
   assign A_pi[0][1][39]  = A_rho[3][0][39];
   assign A_pi[0][1][40]  = A_rho[3][0][40];
   assign A_pi[0][1][41]  = A_rho[3][0][41];
   assign A_pi[0][1][42]  = A_rho[3][0][42];
   assign A_pi[0][1][43]  = A_rho[3][0][43];
   assign A_pi[0][1][44]  = A_rho[3][0][44];
   assign A_pi[0][1][45]  = A_rho[3][0][45];
   assign A_pi[0][1][46]  = A_rho[3][0][46];
   assign A_pi[0][1][47]  = A_rho[3][0][47];
   assign A_pi[0][1][48]  = A_rho[3][0][48];
   assign A_pi[0][1][49]  = A_rho[3][0][49];
   assign A_pi[0][1][50]  = A_rho[3][0][50];
   assign A_pi[0][1][51]  = A_rho[3][0][51];
   assign A_pi[0][1][52]  = A_rho[3][0][52];
   assign A_pi[0][1][53]  = A_rho[3][0][53];
   assign A_pi[0][1][54]  = A_rho[3][0][54];
   assign A_pi[0][1][55]  = A_rho[3][0][55];
   assign A_pi[0][1][56]  = A_rho[3][0][56];
   assign A_pi[0][1][57]  = A_rho[3][0][57];
   assign A_pi[0][1][58]  = A_rho[3][0][58];
   assign A_pi[0][1][59]  = A_rho[3][0][59];
   assign A_pi[0][1][60]  = A_rho[3][0][60];
   assign A_pi[0][1][61]  = A_rho[3][0][61];
   assign A_pi[0][1][62]  = A_rho[3][0][62];
   assign A_pi[0][1][63]  = A_rho[3][0][63];
   assign A_pi[0][2][0]  = A_rho[1][0][0];
   assign A_pi[0][2][1]  = A_rho[1][0][1];
   assign A_pi[0][2][2]  = A_rho[1][0][2];
   assign A_pi[0][2][3]  = A_rho[1][0][3];
   assign A_pi[0][2][4]  = A_rho[1][0][4];
   assign A_pi[0][2][5]  = A_rho[1][0][5];
   assign A_pi[0][2][6]  = A_rho[1][0][6];
   assign A_pi[0][2][7]  = A_rho[1][0][7];
   assign A_pi[0][2][8]  = A_rho[1][0][8];
   assign A_pi[0][2][9]  = A_rho[1][0][9];
   assign A_pi[0][2][10]  = A_rho[1][0][10];
   assign A_pi[0][2][11]  = A_rho[1][0][11];
   assign A_pi[0][2][12]  = A_rho[1][0][12];
   assign A_pi[0][2][13]  = A_rho[1][0][13];
   assign A_pi[0][2][14]  = A_rho[1][0][14];
   assign A_pi[0][2][15]  = A_rho[1][0][15];
   assign A_pi[0][2][16]  = A_rho[1][0][16];
   assign A_pi[0][2][17]  = A_rho[1][0][17];
   assign A_pi[0][2][18]  = A_rho[1][0][18];
   assign A_pi[0][2][19]  = A_rho[1][0][19];
   assign A_pi[0][2][20]  = A_rho[1][0][20];
   assign A_pi[0][2][21]  = A_rho[1][0][21];
   assign A_pi[0][2][22]  = A_rho[1][0][22];
   assign A_pi[0][2][23]  = A_rho[1][0][23];
   assign A_pi[0][2][24]  = A_rho[1][0][24];
   assign A_pi[0][2][25]  = A_rho[1][0][25];
   assign A_pi[0][2][26]  = A_rho[1][0][26];
   assign A_pi[0][2][27]  = A_rho[1][0][27];
   assign A_pi[0][2][28]  = A_rho[1][0][28];
   assign A_pi[0][2][29]  = A_rho[1][0][29];
   assign A_pi[0][2][30]  = A_rho[1][0][30];
   assign A_pi[0][2][31]  = A_rho[1][0][31];
   assign A_pi[0][2][32]  = A_rho[1][0][32];
   assign A_pi[0][2][33]  = A_rho[1][0][33];
   assign A_pi[0][2][34]  = A_rho[1][0][34];
   assign A_pi[0][2][35]  = A_rho[1][0][35];
   assign A_pi[0][2][36]  = A_rho[1][0][36];
   assign A_pi[0][2][37]  = A_rho[1][0][37];
   assign A_pi[0][2][38]  = A_rho[1][0][38];
   assign A_pi[0][2][39]  = A_rho[1][0][39];
   assign A_pi[0][2][40]  = A_rho[1][0][40];
   assign A_pi[0][2][41]  = A_rho[1][0][41];
   assign A_pi[0][2][42]  = A_rho[1][0][42];
   assign A_pi[0][2][43]  = A_rho[1][0][43];
   assign A_pi[0][2][44]  = A_rho[1][0][44];
   assign A_pi[0][2][45]  = A_rho[1][0][45];
   assign A_pi[0][2][46]  = A_rho[1][0][46];
   assign A_pi[0][2][47]  = A_rho[1][0][47];
   assign A_pi[0][2][48]  = A_rho[1][0][48];
   assign A_pi[0][2][49]  = A_rho[1][0][49];
   assign A_pi[0][2][50]  = A_rho[1][0][50];
   assign A_pi[0][2][51]  = A_rho[1][0][51];
   assign A_pi[0][2][52]  = A_rho[1][0][52];
   assign A_pi[0][2][53]  = A_rho[1][0][53];
   assign A_pi[0][2][54]  = A_rho[1][0][54];
   assign A_pi[0][2][55]  = A_rho[1][0][55];
   assign A_pi[0][2][56]  = A_rho[1][0][56];
   assign A_pi[0][2][57]  = A_rho[1][0][57];
   assign A_pi[0][2][58]  = A_rho[1][0][58];
   assign A_pi[0][2][59]  = A_rho[1][0][59];
   assign A_pi[0][2][60]  = A_rho[1][0][60];
   assign A_pi[0][2][61]  = A_rho[1][0][61];
   assign A_pi[0][2][62]  = A_rho[1][0][62];
   assign A_pi[0][2][63]  = A_rho[1][0][63];
   assign A_pi[0][3][0]  = A_rho[4][0][0];
   assign A_pi[0][3][1]  = A_rho[4][0][1];
   assign A_pi[0][3][2]  = A_rho[4][0][2];
   assign A_pi[0][3][3]  = A_rho[4][0][3];
   assign A_pi[0][3][4]  = A_rho[4][0][4];
   assign A_pi[0][3][5]  = A_rho[4][0][5];
   assign A_pi[0][3][6]  = A_rho[4][0][6];
   assign A_pi[0][3][7]  = A_rho[4][0][7];
   assign A_pi[0][3][8]  = A_rho[4][0][8];
   assign A_pi[0][3][9]  = A_rho[4][0][9];
   assign A_pi[0][3][10]  = A_rho[4][0][10];
   assign A_pi[0][3][11]  = A_rho[4][0][11];
   assign A_pi[0][3][12]  = A_rho[4][0][12];
   assign A_pi[0][3][13]  = A_rho[4][0][13];
   assign A_pi[0][3][14]  = A_rho[4][0][14];
   assign A_pi[0][3][15]  = A_rho[4][0][15];
   assign A_pi[0][3][16]  = A_rho[4][0][16];
   assign A_pi[0][3][17]  = A_rho[4][0][17];
   assign A_pi[0][3][18]  = A_rho[4][0][18];
   assign A_pi[0][3][19]  = A_rho[4][0][19];
   assign A_pi[0][3][20]  = A_rho[4][0][20];
   assign A_pi[0][3][21]  = A_rho[4][0][21];
   assign A_pi[0][3][22]  = A_rho[4][0][22];
   assign A_pi[0][3][23]  = A_rho[4][0][23];
   assign A_pi[0][3][24]  = A_rho[4][0][24];
   assign A_pi[0][3][25]  = A_rho[4][0][25];
   assign A_pi[0][3][26]  = A_rho[4][0][26];
   assign A_pi[0][3][27]  = A_rho[4][0][27];
   assign A_pi[0][3][28]  = A_rho[4][0][28];
   assign A_pi[0][3][29]  = A_rho[4][0][29];
   assign A_pi[0][3][30]  = A_rho[4][0][30];
   assign A_pi[0][3][31]  = A_rho[4][0][31];
   assign A_pi[0][3][32]  = A_rho[4][0][32];
   assign A_pi[0][3][33]  = A_rho[4][0][33];
   assign A_pi[0][3][34]  = A_rho[4][0][34];
   assign A_pi[0][3][35]  = A_rho[4][0][35];
   assign A_pi[0][3][36]  = A_rho[4][0][36];
   assign A_pi[0][3][37]  = A_rho[4][0][37];
   assign A_pi[0][3][38]  = A_rho[4][0][38];
   assign A_pi[0][3][39]  = A_rho[4][0][39];
   assign A_pi[0][3][40]  = A_rho[4][0][40];
   assign A_pi[0][3][41]  = A_rho[4][0][41];
   assign A_pi[0][3][42]  = A_rho[4][0][42];
   assign A_pi[0][3][43]  = A_rho[4][0][43];
   assign A_pi[0][3][44]  = A_rho[4][0][44];
   assign A_pi[0][3][45]  = A_rho[4][0][45];
   assign A_pi[0][3][46]  = A_rho[4][0][46];
   assign A_pi[0][3][47]  = A_rho[4][0][47];
   assign A_pi[0][3][48]  = A_rho[4][0][48];
   assign A_pi[0][3][49]  = A_rho[4][0][49];
   assign A_pi[0][3][50]  = A_rho[4][0][50];
   assign A_pi[0][3][51]  = A_rho[4][0][51];
   assign A_pi[0][3][52]  = A_rho[4][0][52];
   assign A_pi[0][3][53]  = A_rho[4][0][53];
   assign A_pi[0][3][54]  = A_rho[4][0][54];
   assign A_pi[0][3][55]  = A_rho[4][0][55];
   assign A_pi[0][3][56]  = A_rho[4][0][56];
   assign A_pi[0][3][57]  = A_rho[4][0][57];
   assign A_pi[0][3][58]  = A_rho[4][0][58];
   assign A_pi[0][3][59]  = A_rho[4][0][59];
   assign A_pi[0][3][60]  = A_rho[4][0][60];
   assign A_pi[0][3][61]  = A_rho[4][0][61];
   assign A_pi[0][3][62]  = A_rho[4][0][62];
   assign A_pi[0][3][63]  = A_rho[4][0][63];
   assign A_pi[0][4][0]  = A_rho[2][0][0];
   assign A_pi[0][4][1]  = A_rho[2][0][1];
   assign A_pi[0][4][2]  = A_rho[2][0][2];
   assign A_pi[0][4][3]  = A_rho[2][0][3];
   assign A_pi[0][4][4]  = A_rho[2][0][4];
   assign A_pi[0][4][5]  = A_rho[2][0][5];
   assign A_pi[0][4][6]  = A_rho[2][0][6];
   assign A_pi[0][4][7]  = A_rho[2][0][7];
   assign A_pi[0][4][8]  = A_rho[2][0][8];
   assign A_pi[0][4][9]  = A_rho[2][0][9];
   assign A_pi[0][4][10]  = A_rho[2][0][10];
   assign A_pi[0][4][11]  = A_rho[2][0][11];
   assign A_pi[0][4][12]  = A_rho[2][0][12];
   assign A_pi[0][4][13]  = A_rho[2][0][13];
   assign A_pi[0][4][14]  = A_rho[2][0][14];
   assign A_pi[0][4][15]  = A_rho[2][0][15];
   assign A_pi[0][4][16]  = A_rho[2][0][16];
   assign A_pi[0][4][17]  = A_rho[2][0][17];
   assign A_pi[0][4][18]  = A_rho[2][0][18];
   assign A_pi[0][4][19]  = A_rho[2][0][19];
   assign A_pi[0][4][20]  = A_rho[2][0][20];
   assign A_pi[0][4][21]  = A_rho[2][0][21];
   assign A_pi[0][4][22]  = A_rho[2][0][22];
   assign A_pi[0][4][23]  = A_rho[2][0][23];
   assign A_pi[0][4][24]  = A_rho[2][0][24];
   assign A_pi[0][4][25]  = A_rho[2][0][25];
   assign A_pi[0][4][26]  = A_rho[2][0][26];
   assign A_pi[0][4][27]  = A_rho[2][0][27];
   assign A_pi[0][4][28]  = A_rho[2][0][28];
   assign A_pi[0][4][29]  = A_rho[2][0][29];
   assign A_pi[0][4][30]  = A_rho[2][0][30];
   assign A_pi[0][4][31]  = A_rho[2][0][31];
   assign A_pi[0][4][32]  = A_rho[2][0][32];
   assign A_pi[0][4][33]  = A_rho[2][0][33];
   assign A_pi[0][4][34]  = A_rho[2][0][34];
   assign A_pi[0][4][35]  = A_rho[2][0][35];
   assign A_pi[0][4][36]  = A_rho[2][0][36];
   assign A_pi[0][4][37]  = A_rho[2][0][37];
   assign A_pi[0][4][38]  = A_rho[2][0][38];
   assign A_pi[0][4][39]  = A_rho[2][0][39];
   assign A_pi[0][4][40]  = A_rho[2][0][40];
   assign A_pi[0][4][41]  = A_rho[2][0][41];
   assign A_pi[0][4][42]  = A_rho[2][0][42];
   assign A_pi[0][4][43]  = A_rho[2][0][43];
   assign A_pi[0][4][44]  = A_rho[2][0][44];
   assign A_pi[0][4][45]  = A_rho[2][0][45];
   assign A_pi[0][4][46]  = A_rho[2][0][46];
   assign A_pi[0][4][47]  = A_rho[2][0][47];
   assign A_pi[0][4][48]  = A_rho[2][0][48];
   assign A_pi[0][4][49]  = A_rho[2][0][49];
   assign A_pi[0][4][50]  = A_rho[2][0][50];
   assign A_pi[0][4][51]  = A_rho[2][0][51];
   assign A_pi[0][4][52]  = A_rho[2][0][52];
   assign A_pi[0][4][53]  = A_rho[2][0][53];
   assign A_pi[0][4][54]  = A_rho[2][0][54];
   assign A_pi[0][4][55]  = A_rho[2][0][55];
   assign A_pi[0][4][56]  = A_rho[2][0][56];
   assign A_pi[0][4][57]  = A_rho[2][0][57];
   assign A_pi[0][4][58]  = A_rho[2][0][58];
   assign A_pi[0][4][59]  = A_rho[2][0][59];
   assign A_pi[0][4][60]  = A_rho[2][0][60];
   assign A_pi[0][4][61]  = A_rho[2][0][61];
   assign A_pi[0][4][62]  = A_rho[2][0][62];
   assign A_pi[0][4][63]  = A_rho[2][0][63];
   assign A_pi[1][0][0]  = A_rho[1][1][0];
   assign A_pi[1][0][1]  = A_rho[1][1][1];
   assign A_pi[1][0][2]  = A_rho[1][1][2];
   assign A_pi[1][0][3]  = A_rho[1][1][3];
   assign A_pi[1][0][4]  = A_rho[1][1][4];
   assign A_pi[1][0][5]  = A_rho[1][1][5];
   assign A_pi[1][0][6]  = A_rho[1][1][6];
   assign A_pi[1][0][7]  = A_rho[1][1][7];
   assign A_pi[1][0][8]  = A_rho[1][1][8];
   assign A_pi[1][0][9]  = A_rho[1][1][9];
   assign A_pi[1][0][10]  = A_rho[1][1][10];
   assign A_pi[1][0][11]  = A_rho[1][1][11];
   assign A_pi[1][0][12]  = A_rho[1][1][12];
   assign A_pi[1][0][13]  = A_rho[1][1][13];
   assign A_pi[1][0][14]  = A_rho[1][1][14];
   assign A_pi[1][0][15]  = A_rho[1][1][15];
   assign A_pi[1][0][16]  = A_rho[1][1][16];
   assign A_pi[1][0][17]  = A_rho[1][1][17];
   assign A_pi[1][0][18]  = A_rho[1][1][18];
   assign A_pi[1][0][19]  = A_rho[1][1][19];
   assign A_pi[1][0][20]  = A_rho[1][1][20];
   assign A_pi[1][0][21]  = A_rho[1][1][21];
   assign A_pi[1][0][22]  = A_rho[1][1][22];
   assign A_pi[1][0][23]  = A_rho[1][1][23];
   assign A_pi[1][0][24]  = A_rho[1][1][24];
   assign A_pi[1][0][25]  = A_rho[1][1][25];
   assign A_pi[1][0][26]  = A_rho[1][1][26];
   assign A_pi[1][0][27]  = A_rho[1][1][27];
   assign A_pi[1][0][28]  = A_rho[1][1][28];
   assign A_pi[1][0][29]  = A_rho[1][1][29];
   assign A_pi[1][0][30]  = A_rho[1][1][30];
   assign A_pi[1][0][31]  = A_rho[1][1][31];
   assign A_pi[1][0][32]  = A_rho[1][1][32];
   assign A_pi[1][0][33]  = A_rho[1][1][33];
   assign A_pi[1][0][34]  = A_rho[1][1][34];
   assign A_pi[1][0][35]  = A_rho[1][1][35];
   assign A_pi[1][0][36]  = A_rho[1][1][36];
   assign A_pi[1][0][37]  = A_rho[1][1][37];
   assign A_pi[1][0][38]  = A_rho[1][1][38];
   assign A_pi[1][0][39]  = A_rho[1][1][39];
   assign A_pi[1][0][40]  = A_rho[1][1][40];
   assign A_pi[1][0][41]  = A_rho[1][1][41];
   assign A_pi[1][0][42]  = A_rho[1][1][42];
   assign A_pi[1][0][43]  = A_rho[1][1][43];
   assign A_pi[1][0][44]  = A_rho[1][1][44];
   assign A_pi[1][0][45]  = A_rho[1][1][45];
   assign A_pi[1][0][46]  = A_rho[1][1][46];
   assign A_pi[1][0][47]  = A_rho[1][1][47];
   assign A_pi[1][0][48]  = A_rho[1][1][48];
   assign A_pi[1][0][49]  = A_rho[1][1][49];
   assign A_pi[1][0][50]  = A_rho[1][1][50];
   assign A_pi[1][0][51]  = A_rho[1][1][51];
   assign A_pi[1][0][52]  = A_rho[1][1][52];
   assign A_pi[1][0][53]  = A_rho[1][1][53];
   assign A_pi[1][0][54]  = A_rho[1][1][54];
   assign A_pi[1][0][55]  = A_rho[1][1][55];
   assign A_pi[1][0][56]  = A_rho[1][1][56];
   assign A_pi[1][0][57]  = A_rho[1][1][57];
   assign A_pi[1][0][58]  = A_rho[1][1][58];
   assign A_pi[1][0][59]  = A_rho[1][1][59];
   assign A_pi[1][0][60]  = A_rho[1][1][60];
   assign A_pi[1][0][61]  = A_rho[1][1][61];
   assign A_pi[1][0][62]  = A_rho[1][1][62];
   assign A_pi[1][0][63]  = A_rho[1][1][63];
   assign A_pi[1][1][0]  = A_rho[4][1][0];
   assign A_pi[1][1][1]  = A_rho[4][1][1];
   assign A_pi[1][1][2]  = A_rho[4][1][2];
   assign A_pi[1][1][3]  = A_rho[4][1][3];
   assign A_pi[1][1][4]  = A_rho[4][1][4];
   assign A_pi[1][1][5]  = A_rho[4][1][5];
   assign A_pi[1][1][6]  = A_rho[4][1][6];
   assign A_pi[1][1][7]  = A_rho[4][1][7];
   assign A_pi[1][1][8]  = A_rho[4][1][8];
   assign A_pi[1][1][9]  = A_rho[4][1][9];
   assign A_pi[1][1][10]  = A_rho[4][1][10];
   assign A_pi[1][1][11]  = A_rho[4][1][11];
   assign A_pi[1][1][12]  = A_rho[4][1][12];
   assign A_pi[1][1][13]  = A_rho[4][1][13];
   assign A_pi[1][1][14]  = A_rho[4][1][14];
   assign A_pi[1][1][15]  = A_rho[4][1][15];
   assign A_pi[1][1][16]  = A_rho[4][1][16];
   assign A_pi[1][1][17]  = A_rho[4][1][17];
   assign A_pi[1][1][18]  = A_rho[4][1][18];
   assign A_pi[1][1][19]  = A_rho[4][1][19];
   assign A_pi[1][1][20]  = A_rho[4][1][20];
   assign A_pi[1][1][21]  = A_rho[4][1][21];
   assign A_pi[1][1][22]  = A_rho[4][1][22];
   assign A_pi[1][1][23]  = A_rho[4][1][23];
   assign A_pi[1][1][24]  = A_rho[4][1][24];
   assign A_pi[1][1][25]  = A_rho[4][1][25];
   assign A_pi[1][1][26]  = A_rho[4][1][26];
   assign A_pi[1][1][27]  = A_rho[4][1][27];
   assign A_pi[1][1][28]  = A_rho[4][1][28];
   assign A_pi[1][1][29]  = A_rho[4][1][29];
   assign A_pi[1][1][30]  = A_rho[4][1][30];
   assign A_pi[1][1][31]  = A_rho[4][1][31];
   assign A_pi[1][1][32]  = A_rho[4][1][32];
   assign A_pi[1][1][33]  = A_rho[4][1][33];
   assign A_pi[1][1][34]  = A_rho[4][1][34];
   assign A_pi[1][1][35]  = A_rho[4][1][35];
   assign A_pi[1][1][36]  = A_rho[4][1][36];
   assign A_pi[1][1][37]  = A_rho[4][1][37];
   assign A_pi[1][1][38]  = A_rho[4][1][38];
   assign A_pi[1][1][39]  = A_rho[4][1][39];
   assign A_pi[1][1][40]  = A_rho[4][1][40];
   assign A_pi[1][1][41]  = A_rho[4][1][41];
   assign A_pi[1][1][42]  = A_rho[4][1][42];
   assign A_pi[1][1][43]  = A_rho[4][1][43];
   assign A_pi[1][1][44]  = A_rho[4][1][44];
   assign A_pi[1][1][45]  = A_rho[4][1][45];
   assign A_pi[1][1][46]  = A_rho[4][1][46];
   assign A_pi[1][1][47]  = A_rho[4][1][47];
   assign A_pi[1][1][48]  = A_rho[4][1][48];
   assign A_pi[1][1][49]  = A_rho[4][1][49];
   assign A_pi[1][1][50]  = A_rho[4][1][50];
   assign A_pi[1][1][51]  = A_rho[4][1][51];
   assign A_pi[1][1][52]  = A_rho[4][1][52];
   assign A_pi[1][1][53]  = A_rho[4][1][53];
   assign A_pi[1][1][54]  = A_rho[4][1][54];
   assign A_pi[1][1][55]  = A_rho[4][1][55];
   assign A_pi[1][1][56]  = A_rho[4][1][56];
   assign A_pi[1][1][57]  = A_rho[4][1][57];
   assign A_pi[1][1][58]  = A_rho[4][1][58];
   assign A_pi[1][1][59]  = A_rho[4][1][59];
   assign A_pi[1][1][60]  = A_rho[4][1][60];
   assign A_pi[1][1][61]  = A_rho[4][1][61];
   assign A_pi[1][1][62]  = A_rho[4][1][62];
   assign A_pi[1][1][63]  = A_rho[4][1][63];
   assign A_pi[1][2][0]  = A_rho[2][1][0];
   assign A_pi[1][2][1]  = A_rho[2][1][1];
   assign A_pi[1][2][2]  = A_rho[2][1][2];
   assign A_pi[1][2][3]  = A_rho[2][1][3];
   assign A_pi[1][2][4]  = A_rho[2][1][4];
   assign A_pi[1][2][5]  = A_rho[2][1][5];
   assign A_pi[1][2][6]  = A_rho[2][1][6];
   assign A_pi[1][2][7]  = A_rho[2][1][7];
   assign A_pi[1][2][8]  = A_rho[2][1][8];
   assign A_pi[1][2][9]  = A_rho[2][1][9];
   assign A_pi[1][2][10]  = A_rho[2][1][10];
   assign A_pi[1][2][11]  = A_rho[2][1][11];
   assign A_pi[1][2][12]  = A_rho[2][1][12];
   assign A_pi[1][2][13]  = A_rho[2][1][13];
   assign A_pi[1][2][14]  = A_rho[2][1][14];
   assign A_pi[1][2][15]  = A_rho[2][1][15];
   assign A_pi[1][2][16]  = A_rho[2][1][16];
   assign A_pi[1][2][17]  = A_rho[2][1][17];
   assign A_pi[1][2][18]  = A_rho[2][1][18];
   assign A_pi[1][2][19]  = A_rho[2][1][19];
   assign A_pi[1][2][20]  = A_rho[2][1][20];
   assign A_pi[1][2][21]  = A_rho[2][1][21];
   assign A_pi[1][2][22]  = A_rho[2][1][22];
   assign A_pi[1][2][23]  = A_rho[2][1][23];
   assign A_pi[1][2][24]  = A_rho[2][1][24];
   assign A_pi[1][2][25]  = A_rho[2][1][25];
   assign A_pi[1][2][26]  = A_rho[2][1][26];
   assign A_pi[1][2][27]  = A_rho[2][1][27];
   assign A_pi[1][2][28]  = A_rho[2][1][28];
   assign A_pi[1][2][29]  = A_rho[2][1][29];
   assign A_pi[1][2][30]  = A_rho[2][1][30];
   assign A_pi[1][2][31]  = A_rho[2][1][31];
   assign A_pi[1][2][32]  = A_rho[2][1][32];
   assign A_pi[1][2][33]  = A_rho[2][1][33];
   assign A_pi[1][2][34]  = A_rho[2][1][34];
   assign A_pi[1][2][35]  = A_rho[2][1][35];
   assign A_pi[1][2][36]  = A_rho[2][1][36];
   assign A_pi[1][2][37]  = A_rho[2][1][37];
   assign A_pi[1][2][38]  = A_rho[2][1][38];
   assign A_pi[1][2][39]  = A_rho[2][1][39];
   assign A_pi[1][2][40]  = A_rho[2][1][40];
   assign A_pi[1][2][41]  = A_rho[2][1][41];
   assign A_pi[1][2][42]  = A_rho[2][1][42];
   assign A_pi[1][2][43]  = A_rho[2][1][43];
   assign A_pi[1][2][44]  = A_rho[2][1][44];
   assign A_pi[1][2][45]  = A_rho[2][1][45];
   assign A_pi[1][2][46]  = A_rho[2][1][46];
   assign A_pi[1][2][47]  = A_rho[2][1][47];
   assign A_pi[1][2][48]  = A_rho[2][1][48];
   assign A_pi[1][2][49]  = A_rho[2][1][49];
   assign A_pi[1][2][50]  = A_rho[2][1][50];
   assign A_pi[1][2][51]  = A_rho[2][1][51];
   assign A_pi[1][2][52]  = A_rho[2][1][52];
   assign A_pi[1][2][53]  = A_rho[2][1][53];
   assign A_pi[1][2][54]  = A_rho[2][1][54];
   assign A_pi[1][2][55]  = A_rho[2][1][55];
   assign A_pi[1][2][56]  = A_rho[2][1][56];
   assign A_pi[1][2][57]  = A_rho[2][1][57];
   assign A_pi[1][2][58]  = A_rho[2][1][58];
   assign A_pi[1][2][59]  = A_rho[2][1][59];
   assign A_pi[1][2][60]  = A_rho[2][1][60];
   assign A_pi[1][2][61]  = A_rho[2][1][61];
   assign A_pi[1][2][62]  = A_rho[2][1][62];
   assign A_pi[1][2][63]  = A_rho[2][1][63];
   assign A_pi[1][3][0]  = A_rho[0][1][0];
   assign A_pi[1][3][1]  = A_rho[0][1][1];
   assign A_pi[1][3][2]  = A_rho[0][1][2];
   assign A_pi[1][3][3]  = A_rho[0][1][3];
   assign A_pi[1][3][4]  = A_rho[0][1][4];
   assign A_pi[1][3][5]  = A_rho[0][1][5];
   assign A_pi[1][3][6]  = A_rho[0][1][6];
   assign A_pi[1][3][7]  = A_rho[0][1][7];
   assign A_pi[1][3][8]  = A_rho[0][1][8];
   assign A_pi[1][3][9]  = A_rho[0][1][9];
   assign A_pi[1][3][10]  = A_rho[0][1][10];
   assign A_pi[1][3][11]  = A_rho[0][1][11];
   assign A_pi[1][3][12]  = A_rho[0][1][12];
   assign A_pi[1][3][13]  = A_rho[0][1][13];
   assign A_pi[1][3][14]  = A_rho[0][1][14];
   assign A_pi[1][3][15]  = A_rho[0][1][15];
   assign A_pi[1][3][16]  = A_rho[0][1][16];
   assign A_pi[1][3][17]  = A_rho[0][1][17];
   assign A_pi[1][3][18]  = A_rho[0][1][18];
   assign A_pi[1][3][19]  = A_rho[0][1][19];
   assign A_pi[1][3][20]  = A_rho[0][1][20];
   assign A_pi[1][3][21]  = A_rho[0][1][21];
   assign A_pi[1][3][22]  = A_rho[0][1][22];
   assign A_pi[1][3][23]  = A_rho[0][1][23];
   assign A_pi[1][3][24]  = A_rho[0][1][24];
   assign A_pi[1][3][25]  = A_rho[0][1][25];
   assign A_pi[1][3][26]  = A_rho[0][1][26];
   assign A_pi[1][3][27]  = A_rho[0][1][27];
   assign A_pi[1][3][28]  = A_rho[0][1][28];
   assign A_pi[1][3][29]  = A_rho[0][1][29];
   assign A_pi[1][3][30]  = A_rho[0][1][30];
   assign A_pi[1][3][31]  = A_rho[0][1][31];
   assign A_pi[1][3][32]  = A_rho[0][1][32];
   assign A_pi[1][3][33]  = A_rho[0][1][33];
   assign A_pi[1][3][34]  = A_rho[0][1][34];
   assign A_pi[1][3][35]  = A_rho[0][1][35];
   assign A_pi[1][3][36]  = A_rho[0][1][36];
   assign A_pi[1][3][37]  = A_rho[0][1][37];
   assign A_pi[1][3][38]  = A_rho[0][1][38];
   assign A_pi[1][3][39]  = A_rho[0][1][39];
   assign A_pi[1][3][40]  = A_rho[0][1][40];
   assign A_pi[1][3][41]  = A_rho[0][1][41];
   assign A_pi[1][3][42]  = A_rho[0][1][42];
   assign A_pi[1][3][43]  = A_rho[0][1][43];
   assign A_pi[1][3][44]  = A_rho[0][1][44];
   assign A_pi[1][3][45]  = A_rho[0][1][45];
   assign A_pi[1][3][46]  = A_rho[0][1][46];
   assign A_pi[1][3][47]  = A_rho[0][1][47];
   assign A_pi[1][3][48]  = A_rho[0][1][48];
   assign A_pi[1][3][49]  = A_rho[0][1][49];
   assign A_pi[1][3][50]  = A_rho[0][1][50];
   assign A_pi[1][3][51]  = A_rho[0][1][51];
   assign A_pi[1][3][52]  = A_rho[0][1][52];
   assign A_pi[1][3][53]  = A_rho[0][1][53];
   assign A_pi[1][3][54]  = A_rho[0][1][54];
   assign A_pi[1][3][55]  = A_rho[0][1][55];
   assign A_pi[1][3][56]  = A_rho[0][1][56];
   assign A_pi[1][3][57]  = A_rho[0][1][57];
   assign A_pi[1][3][58]  = A_rho[0][1][58];
   assign A_pi[1][3][59]  = A_rho[0][1][59];
   assign A_pi[1][3][60]  = A_rho[0][1][60];
   assign A_pi[1][3][61]  = A_rho[0][1][61];
   assign A_pi[1][3][62]  = A_rho[0][1][62];
   assign A_pi[1][3][63]  = A_rho[0][1][63];
   assign A_pi[1][4][0]  = A_rho[3][1][0];
   assign A_pi[1][4][1]  = A_rho[3][1][1];
   assign A_pi[1][4][2]  = A_rho[3][1][2];
   assign A_pi[1][4][3]  = A_rho[3][1][3];
   assign A_pi[1][4][4]  = A_rho[3][1][4];
   assign A_pi[1][4][5]  = A_rho[3][1][5];
   assign A_pi[1][4][6]  = A_rho[3][1][6];
   assign A_pi[1][4][7]  = A_rho[3][1][7];
   assign A_pi[1][4][8]  = A_rho[3][1][8];
   assign A_pi[1][4][9]  = A_rho[3][1][9];
   assign A_pi[1][4][10]  = A_rho[3][1][10];
   assign A_pi[1][4][11]  = A_rho[3][1][11];
   assign A_pi[1][4][12]  = A_rho[3][1][12];
   assign A_pi[1][4][13]  = A_rho[3][1][13];
   assign A_pi[1][4][14]  = A_rho[3][1][14];
   assign A_pi[1][4][15]  = A_rho[3][1][15];
   assign A_pi[1][4][16]  = A_rho[3][1][16];
   assign A_pi[1][4][17]  = A_rho[3][1][17];
   assign A_pi[1][4][18]  = A_rho[3][1][18];
   assign A_pi[1][4][19]  = A_rho[3][1][19];
   assign A_pi[1][4][20]  = A_rho[3][1][20];
   assign A_pi[1][4][21]  = A_rho[3][1][21];
   assign A_pi[1][4][22]  = A_rho[3][1][22];
   assign A_pi[1][4][23]  = A_rho[3][1][23];
   assign A_pi[1][4][24]  = A_rho[3][1][24];
   assign A_pi[1][4][25]  = A_rho[3][1][25];
   assign A_pi[1][4][26]  = A_rho[3][1][26];
   assign A_pi[1][4][27]  = A_rho[3][1][27];
   assign A_pi[1][4][28]  = A_rho[3][1][28];
   assign A_pi[1][4][29]  = A_rho[3][1][29];
   assign A_pi[1][4][30]  = A_rho[3][1][30];
   assign A_pi[1][4][31]  = A_rho[3][1][31];
   assign A_pi[1][4][32]  = A_rho[3][1][32];
   assign A_pi[1][4][33]  = A_rho[3][1][33];
   assign A_pi[1][4][34]  = A_rho[3][1][34];
   assign A_pi[1][4][35]  = A_rho[3][1][35];
   assign A_pi[1][4][36]  = A_rho[3][1][36];
   assign A_pi[1][4][37]  = A_rho[3][1][37];
   assign A_pi[1][4][38]  = A_rho[3][1][38];
   assign A_pi[1][4][39]  = A_rho[3][1][39];
   assign A_pi[1][4][40]  = A_rho[3][1][40];
   assign A_pi[1][4][41]  = A_rho[3][1][41];
   assign A_pi[1][4][42]  = A_rho[3][1][42];
   assign A_pi[1][4][43]  = A_rho[3][1][43];
   assign A_pi[1][4][44]  = A_rho[3][1][44];
   assign A_pi[1][4][45]  = A_rho[3][1][45];
   assign A_pi[1][4][46]  = A_rho[3][1][46];
   assign A_pi[1][4][47]  = A_rho[3][1][47];
   assign A_pi[1][4][48]  = A_rho[3][1][48];
   assign A_pi[1][4][49]  = A_rho[3][1][49];
   assign A_pi[1][4][50]  = A_rho[3][1][50];
   assign A_pi[1][4][51]  = A_rho[3][1][51];
   assign A_pi[1][4][52]  = A_rho[3][1][52];
   assign A_pi[1][4][53]  = A_rho[3][1][53];
   assign A_pi[1][4][54]  = A_rho[3][1][54];
   assign A_pi[1][4][55]  = A_rho[3][1][55];
   assign A_pi[1][4][56]  = A_rho[3][1][56];
   assign A_pi[1][4][57]  = A_rho[3][1][57];
   assign A_pi[1][4][58]  = A_rho[3][1][58];
   assign A_pi[1][4][59]  = A_rho[3][1][59];
   assign A_pi[1][4][60]  = A_rho[3][1][60];
   assign A_pi[1][4][61]  = A_rho[3][1][61];
   assign A_pi[1][4][62]  = A_rho[3][1][62];
   assign A_pi[1][4][63]  = A_rho[3][1][63];
   assign A_pi[2][0][0]  = A_rho[2][2][0];
   assign A_pi[2][0][1]  = A_rho[2][2][1];
   assign A_pi[2][0][2]  = A_rho[2][2][2];
   assign A_pi[2][0][3]  = A_rho[2][2][3];
   assign A_pi[2][0][4]  = A_rho[2][2][4];
   assign A_pi[2][0][5]  = A_rho[2][2][5];
   assign A_pi[2][0][6]  = A_rho[2][2][6];
   assign A_pi[2][0][7]  = A_rho[2][2][7];
   assign A_pi[2][0][8]  = A_rho[2][2][8];
   assign A_pi[2][0][9]  = A_rho[2][2][9];
   assign A_pi[2][0][10]  = A_rho[2][2][10];
   assign A_pi[2][0][11]  = A_rho[2][2][11];
   assign A_pi[2][0][12]  = A_rho[2][2][12];
   assign A_pi[2][0][13]  = A_rho[2][2][13];
   assign A_pi[2][0][14]  = A_rho[2][2][14];
   assign A_pi[2][0][15]  = A_rho[2][2][15];
   assign A_pi[2][0][16]  = A_rho[2][2][16];
   assign A_pi[2][0][17]  = A_rho[2][2][17];
   assign A_pi[2][0][18]  = A_rho[2][2][18];
   assign A_pi[2][0][19]  = A_rho[2][2][19];
   assign A_pi[2][0][20]  = A_rho[2][2][20];
   assign A_pi[2][0][21]  = A_rho[2][2][21];
   assign A_pi[2][0][22]  = A_rho[2][2][22];
   assign A_pi[2][0][23]  = A_rho[2][2][23];
   assign A_pi[2][0][24]  = A_rho[2][2][24];
   assign A_pi[2][0][25]  = A_rho[2][2][25];
   assign A_pi[2][0][26]  = A_rho[2][2][26];
   assign A_pi[2][0][27]  = A_rho[2][2][27];
   assign A_pi[2][0][28]  = A_rho[2][2][28];
   assign A_pi[2][0][29]  = A_rho[2][2][29];
   assign A_pi[2][0][30]  = A_rho[2][2][30];
   assign A_pi[2][0][31]  = A_rho[2][2][31];
   assign A_pi[2][0][32]  = A_rho[2][2][32];
   assign A_pi[2][0][33]  = A_rho[2][2][33];
   assign A_pi[2][0][34]  = A_rho[2][2][34];
   assign A_pi[2][0][35]  = A_rho[2][2][35];
   assign A_pi[2][0][36]  = A_rho[2][2][36];
   assign A_pi[2][0][37]  = A_rho[2][2][37];
   assign A_pi[2][0][38]  = A_rho[2][2][38];
   assign A_pi[2][0][39]  = A_rho[2][2][39];
   assign A_pi[2][0][40]  = A_rho[2][2][40];
   assign A_pi[2][0][41]  = A_rho[2][2][41];
   assign A_pi[2][0][42]  = A_rho[2][2][42];
   assign A_pi[2][0][43]  = A_rho[2][2][43];
   assign A_pi[2][0][44]  = A_rho[2][2][44];
   assign A_pi[2][0][45]  = A_rho[2][2][45];
   assign A_pi[2][0][46]  = A_rho[2][2][46];
   assign A_pi[2][0][47]  = A_rho[2][2][47];
   assign A_pi[2][0][48]  = A_rho[2][2][48];
   assign A_pi[2][0][49]  = A_rho[2][2][49];
   assign A_pi[2][0][50]  = A_rho[2][2][50];
   assign A_pi[2][0][51]  = A_rho[2][2][51];
   assign A_pi[2][0][52]  = A_rho[2][2][52];
   assign A_pi[2][0][53]  = A_rho[2][2][53];
   assign A_pi[2][0][54]  = A_rho[2][2][54];
   assign A_pi[2][0][55]  = A_rho[2][2][55];
   assign A_pi[2][0][56]  = A_rho[2][2][56];
   assign A_pi[2][0][57]  = A_rho[2][2][57];
   assign A_pi[2][0][58]  = A_rho[2][2][58];
   assign A_pi[2][0][59]  = A_rho[2][2][59];
   assign A_pi[2][0][60]  = A_rho[2][2][60];
   assign A_pi[2][0][61]  = A_rho[2][2][61];
   assign A_pi[2][0][62]  = A_rho[2][2][62];
   assign A_pi[2][0][63]  = A_rho[2][2][63];
   assign A_pi[2][1][0]  = A_rho[0][2][0];
   assign A_pi[2][1][1]  = A_rho[0][2][1];
   assign A_pi[2][1][2]  = A_rho[0][2][2];
   assign A_pi[2][1][3]  = A_rho[0][2][3];
   assign A_pi[2][1][4]  = A_rho[0][2][4];
   assign A_pi[2][1][5]  = A_rho[0][2][5];
   assign A_pi[2][1][6]  = A_rho[0][2][6];
   assign A_pi[2][1][7]  = A_rho[0][2][7];
   assign A_pi[2][1][8]  = A_rho[0][2][8];
   assign A_pi[2][1][9]  = A_rho[0][2][9];
   assign A_pi[2][1][10]  = A_rho[0][2][10];
   assign A_pi[2][1][11]  = A_rho[0][2][11];
   assign A_pi[2][1][12]  = A_rho[0][2][12];
   assign A_pi[2][1][13]  = A_rho[0][2][13];
   assign A_pi[2][1][14]  = A_rho[0][2][14];
   assign A_pi[2][1][15]  = A_rho[0][2][15];
   assign A_pi[2][1][16]  = A_rho[0][2][16];
   assign A_pi[2][1][17]  = A_rho[0][2][17];
   assign A_pi[2][1][18]  = A_rho[0][2][18];
   assign A_pi[2][1][19]  = A_rho[0][2][19];
   assign A_pi[2][1][20]  = A_rho[0][2][20];
   assign A_pi[2][1][21]  = A_rho[0][2][21];
   assign A_pi[2][1][22]  = A_rho[0][2][22];
   assign A_pi[2][1][23]  = A_rho[0][2][23];
   assign A_pi[2][1][24]  = A_rho[0][2][24];
   assign A_pi[2][1][25]  = A_rho[0][2][25];
   assign A_pi[2][1][26]  = A_rho[0][2][26];
   assign A_pi[2][1][27]  = A_rho[0][2][27];
   assign A_pi[2][1][28]  = A_rho[0][2][28];
   assign A_pi[2][1][29]  = A_rho[0][2][29];
   assign A_pi[2][1][30]  = A_rho[0][2][30];
   assign A_pi[2][1][31]  = A_rho[0][2][31];
   assign A_pi[2][1][32]  = A_rho[0][2][32];
   assign A_pi[2][1][33]  = A_rho[0][2][33];
   assign A_pi[2][1][34]  = A_rho[0][2][34];
   assign A_pi[2][1][35]  = A_rho[0][2][35];
   assign A_pi[2][1][36]  = A_rho[0][2][36];
   assign A_pi[2][1][37]  = A_rho[0][2][37];
   assign A_pi[2][1][38]  = A_rho[0][2][38];
   assign A_pi[2][1][39]  = A_rho[0][2][39];
   assign A_pi[2][1][40]  = A_rho[0][2][40];
   assign A_pi[2][1][41]  = A_rho[0][2][41];
   assign A_pi[2][1][42]  = A_rho[0][2][42];
   assign A_pi[2][1][43]  = A_rho[0][2][43];
   assign A_pi[2][1][44]  = A_rho[0][2][44];
   assign A_pi[2][1][45]  = A_rho[0][2][45];
   assign A_pi[2][1][46]  = A_rho[0][2][46];
   assign A_pi[2][1][47]  = A_rho[0][2][47];
   assign A_pi[2][1][48]  = A_rho[0][2][48];
   assign A_pi[2][1][49]  = A_rho[0][2][49];
   assign A_pi[2][1][50]  = A_rho[0][2][50];
   assign A_pi[2][1][51]  = A_rho[0][2][51];
   assign A_pi[2][1][52]  = A_rho[0][2][52];
   assign A_pi[2][1][53]  = A_rho[0][2][53];
   assign A_pi[2][1][54]  = A_rho[0][2][54];
   assign A_pi[2][1][55]  = A_rho[0][2][55];
   assign A_pi[2][1][56]  = A_rho[0][2][56];
   assign A_pi[2][1][57]  = A_rho[0][2][57];
   assign A_pi[2][1][58]  = A_rho[0][2][58];
   assign A_pi[2][1][59]  = A_rho[0][2][59];
   assign A_pi[2][1][60]  = A_rho[0][2][60];
   assign A_pi[2][1][61]  = A_rho[0][2][61];
   assign A_pi[2][1][62]  = A_rho[0][2][62];
   assign A_pi[2][1][63]  = A_rho[0][2][63];
   assign A_pi[2][2][0]  = A_rho[3][2][0];
   assign A_pi[2][2][1]  = A_rho[3][2][1];
   assign A_pi[2][2][2]  = A_rho[3][2][2];
   assign A_pi[2][2][3]  = A_rho[3][2][3];
   assign A_pi[2][2][4]  = A_rho[3][2][4];
   assign A_pi[2][2][5]  = A_rho[3][2][5];
   assign A_pi[2][2][6]  = A_rho[3][2][6];
   assign A_pi[2][2][7]  = A_rho[3][2][7];
   assign A_pi[2][2][8]  = A_rho[3][2][8];
   assign A_pi[2][2][9]  = A_rho[3][2][9];
   assign A_pi[2][2][10]  = A_rho[3][2][10];
   assign A_pi[2][2][11]  = A_rho[3][2][11];
   assign A_pi[2][2][12]  = A_rho[3][2][12];
   assign A_pi[2][2][13]  = A_rho[3][2][13];
   assign A_pi[2][2][14]  = A_rho[3][2][14];
   assign A_pi[2][2][15]  = A_rho[3][2][15];
   assign A_pi[2][2][16]  = A_rho[3][2][16];
   assign A_pi[2][2][17]  = A_rho[3][2][17];
   assign A_pi[2][2][18]  = A_rho[3][2][18];
   assign A_pi[2][2][19]  = A_rho[3][2][19];
   assign A_pi[2][2][20]  = A_rho[3][2][20];
   assign A_pi[2][2][21]  = A_rho[3][2][21];
   assign A_pi[2][2][22]  = A_rho[3][2][22];
   assign A_pi[2][2][23]  = A_rho[3][2][23];
   assign A_pi[2][2][24]  = A_rho[3][2][24];
   assign A_pi[2][2][25]  = A_rho[3][2][25];
   assign A_pi[2][2][26]  = A_rho[3][2][26];
   assign A_pi[2][2][27]  = A_rho[3][2][27];
   assign A_pi[2][2][28]  = A_rho[3][2][28];
   assign A_pi[2][2][29]  = A_rho[3][2][29];
   assign A_pi[2][2][30]  = A_rho[3][2][30];
   assign A_pi[2][2][31]  = A_rho[3][2][31];
   assign A_pi[2][2][32]  = A_rho[3][2][32];
   assign A_pi[2][2][33]  = A_rho[3][2][33];
   assign A_pi[2][2][34]  = A_rho[3][2][34];
   assign A_pi[2][2][35]  = A_rho[3][2][35];
   assign A_pi[2][2][36]  = A_rho[3][2][36];
   assign A_pi[2][2][37]  = A_rho[3][2][37];
   assign A_pi[2][2][38]  = A_rho[3][2][38];
   assign A_pi[2][2][39]  = A_rho[3][2][39];
   assign A_pi[2][2][40]  = A_rho[3][2][40];
   assign A_pi[2][2][41]  = A_rho[3][2][41];
   assign A_pi[2][2][42]  = A_rho[3][2][42];
   assign A_pi[2][2][43]  = A_rho[3][2][43];
   assign A_pi[2][2][44]  = A_rho[3][2][44];
   assign A_pi[2][2][45]  = A_rho[3][2][45];
   assign A_pi[2][2][46]  = A_rho[3][2][46];
   assign A_pi[2][2][47]  = A_rho[3][2][47];
   assign A_pi[2][2][48]  = A_rho[3][2][48];
   assign A_pi[2][2][49]  = A_rho[3][2][49];
   assign A_pi[2][2][50]  = A_rho[3][2][50];
   assign A_pi[2][2][51]  = A_rho[3][2][51];
   assign A_pi[2][2][52]  = A_rho[3][2][52];
   assign A_pi[2][2][53]  = A_rho[3][2][53];
   assign A_pi[2][2][54]  = A_rho[3][2][54];
   assign A_pi[2][2][55]  = A_rho[3][2][55];
   assign A_pi[2][2][56]  = A_rho[3][2][56];
   assign A_pi[2][2][57]  = A_rho[3][2][57];
   assign A_pi[2][2][58]  = A_rho[3][2][58];
   assign A_pi[2][2][59]  = A_rho[3][2][59];
   assign A_pi[2][2][60]  = A_rho[3][2][60];
   assign A_pi[2][2][61]  = A_rho[3][2][61];
   assign A_pi[2][2][62]  = A_rho[3][2][62];
   assign A_pi[2][2][63]  = A_rho[3][2][63];
   assign A_pi[2][3][0]  = A_rho[1][2][0];
   assign A_pi[2][3][1]  = A_rho[1][2][1];
   assign A_pi[2][3][2]  = A_rho[1][2][2];
   assign A_pi[2][3][3]  = A_rho[1][2][3];
   assign A_pi[2][3][4]  = A_rho[1][2][4];
   assign A_pi[2][3][5]  = A_rho[1][2][5];
   assign A_pi[2][3][6]  = A_rho[1][2][6];
   assign A_pi[2][3][7]  = A_rho[1][2][7];
   assign A_pi[2][3][8]  = A_rho[1][2][8];
   assign A_pi[2][3][9]  = A_rho[1][2][9];
   assign A_pi[2][3][10]  = A_rho[1][2][10];
   assign A_pi[2][3][11]  = A_rho[1][2][11];
   assign A_pi[2][3][12]  = A_rho[1][2][12];
   assign A_pi[2][3][13]  = A_rho[1][2][13];
   assign A_pi[2][3][14]  = A_rho[1][2][14];
   assign A_pi[2][3][15]  = A_rho[1][2][15];
   assign A_pi[2][3][16]  = A_rho[1][2][16];
   assign A_pi[2][3][17]  = A_rho[1][2][17];
   assign A_pi[2][3][18]  = A_rho[1][2][18];
   assign A_pi[2][3][19]  = A_rho[1][2][19];
   assign A_pi[2][3][20]  = A_rho[1][2][20];
   assign A_pi[2][3][21]  = A_rho[1][2][21];
   assign A_pi[2][3][22]  = A_rho[1][2][22];
   assign A_pi[2][3][23]  = A_rho[1][2][23];
   assign A_pi[2][3][24]  = A_rho[1][2][24];
   assign A_pi[2][3][25]  = A_rho[1][2][25];
   assign A_pi[2][3][26]  = A_rho[1][2][26];
   assign A_pi[2][3][27]  = A_rho[1][2][27];
   assign A_pi[2][3][28]  = A_rho[1][2][28];
   assign A_pi[2][3][29]  = A_rho[1][2][29];
   assign A_pi[2][3][30]  = A_rho[1][2][30];
   assign A_pi[2][3][31]  = A_rho[1][2][31];
   assign A_pi[2][3][32]  = A_rho[1][2][32];
   assign A_pi[2][3][33]  = A_rho[1][2][33];
   assign A_pi[2][3][34]  = A_rho[1][2][34];
   assign A_pi[2][3][35]  = A_rho[1][2][35];
   assign A_pi[2][3][36]  = A_rho[1][2][36];
   assign A_pi[2][3][37]  = A_rho[1][2][37];
   assign A_pi[2][3][38]  = A_rho[1][2][38];
   assign A_pi[2][3][39]  = A_rho[1][2][39];
   assign A_pi[2][3][40]  = A_rho[1][2][40];
   assign A_pi[2][3][41]  = A_rho[1][2][41];
   assign A_pi[2][3][42]  = A_rho[1][2][42];
   assign A_pi[2][3][43]  = A_rho[1][2][43];
   assign A_pi[2][3][44]  = A_rho[1][2][44];
   assign A_pi[2][3][45]  = A_rho[1][2][45];
   assign A_pi[2][3][46]  = A_rho[1][2][46];
   assign A_pi[2][3][47]  = A_rho[1][2][47];
   assign A_pi[2][3][48]  = A_rho[1][2][48];
   assign A_pi[2][3][49]  = A_rho[1][2][49];
   assign A_pi[2][3][50]  = A_rho[1][2][50];
   assign A_pi[2][3][51]  = A_rho[1][2][51];
   assign A_pi[2][3][52]  = A_rho[1][2][52];
   assign A_pi[2][3][53]  = A_rho[1][2][53];
   assign A_pi[2][3][54]  = A_rho[1][2][54];
   assign A_pi[2][3][55]  = A_rho[1][2][55];
   assign A_pi[2][3][56]  = A_rho[1][2][56];
   assign A_pi[2][3][57]  = A_rho[1][2][57];
   assign A_pi[2][3][58]  = A_rho[1][2][58];
   assign A_pi[2][3][59]  = A_rho[1][2][59];
   assign A_pi[2][3][60]  = A_rho[1][2][60];
   assign A_pi[2][3][61]  = A_rho[1][2][61];
   assign A_pi[2][3][62]  = A_rho[1][2][62];
   assign A_pi[2][3][63]  = A_rho[1][2][63];
   assign A_pi[2][4][0]  = A_rho[4][2][0];
   assign A_pi[2][4][1]  = A_rho[4][2][1];
   assign A_pi[2][4][2]  = A_rho[4][2][2];
   assign A_pi[2][4][3]  = A_rho[4][2][3];
   assign A_pi[2][4][4]  = A_rho[4][2][4];
   assign A_pi[2][4][5]  = A_rho[4][2][5];
   assign A_pi[2][4][6]  = A_rho[4][2][6];
   assign A_pi[2][4][7]  = A_rho[4][2][7];
   assign A_pi[2][4][8]  = A_rho[4][2][8];
   assign A_pi[2][4][9]  = A_rho[4][2][9];
   assign A_pi[2][4][10]  = A_rho[4][2][10];
   assign A_pi[2][4][11]  = A_rho[4][2][11];
   assign A_pi[2][4][12]  = A_rho[4][2][12];
   assign A_pi[2][4][13]  = A_rho[4][2][13];
   assign A_pi[2][4][14]  = A_rho[4][2][14];
   assign A_pi[2][4][15]  = A_rho[4][2][15];
   assign A_pi[2][4][16]  = A_rho[4][2][16];
   assign A_pi[2][4][17]  = A_rho[4][2][17];
   assign A_pi[2][4][18]  = A_rho[4][2][18];
   assign A_pi[2][4][19]  = A_rho[4][2][19];
   assign A_pi[2][4][20]  = A_rho[4][2][20];
   assign A_pi[2][4][21]  = A_rho[4][2][21];
   assign A_pi[2][4][22]  = A_rho[4][2][22];
   assign A_pi[2][4][23]  = A_rho[4][2][23];
   assign A_pi[2][4][24]  = A_rho[4][2][24];
   assign A_pi[2][4][25]  = A_rho[4][2][25];
   assign A_pi[2][4][26]  = A_rho[4][2][26];
   assign A_pi[2][4][27]  = A_rho[4][2][27];
   assign A_pi[2][4][28]  = A_rho[4][2][28];
   assign A_pi[2][4][29]  = A_rho[4][2][29];
   assign A_pi[2][4][30]  = A_rho[4][2][30];
   assign A_pi[2][4][31]  = A_rho[4][2][31];
   assign A_pi[2][4][32]  = A_rho[4][2][32];
   assign A_pi[2][4][33]  = A_rho[4][2][33];
   assign A_pi[2][4][34]  = A_rho[4][2][34];
   assign A_pi[2][4][35]  = A_rho[4][2][35];
   assign A_pi[2][4][36]  = A_rho[4][2][36];
   assign A_pi[2][4][37]  = A_rho[4][2][37];
   assign A_pi[2][4][38]  = A_rho[4][2][38];
   assign A_pi[2][4][39]  = A_rho[4][2][39];
   assign A_pi[2][4][40]  = A_rho[4][2][40];
   assign A_pi[2][4][41]  = A_rho[4][2][41];
   assign A_pi[2][4][42]  = A_rho[4][2][42];
   assign A_pi[2][4][43]  = A_rho[4][2][43];
   assign A_pi[2][4][44]  = A_rho[4][2][44];
   assign A_pi[2][4][45]  = A_rho[4][2][45];
   assign A_pi[2][4][46]  = A_rho[4][2][46];
   assign A_pi[2][4][47]  = A_rho[4][2][47];
   assign A_pi[2][4][48]  = A_rho[4][2][48];
   assign A_pi[2][4][49]  = A_rho[4][2][49];
   assign A_pi[2][4][50]  = A_rho[4][2][50];
   assign A_pi[2][4][51]  = A_rho[4][2][51];
   assign A_pi[2][4][52]  = A_rho[4][2][52];
   assign A_pi[2][4][53]  = A_rho[4][2][53];
   assign A_pi[2][4][54]  = A_rho[4][2][54];
   assign A_pi[2][4][55]  = A_rho[4][2][55];
   assign A_pi[2][4][56]  = A_rho[4][2][56];
   assign A_pi[2][4][57]  = A_rho[4][2][57];
   assign A_pi[2][4][58]  = A_rho[4][2][58];
   assign A_pi[2][4][59]  = A_rho[4][2][59];
   assign A_pi[2][4][60]  = A_rho[4][2][60];
   assign A_pi[2][4][61]  = A_rho[4][2][61];
   assign A_pi[2][4][62]  = A_rho[4][2][62];
   assign A_pi[2][4][63]  = A_rho[4][2][63];
   assign A_pi[3][0][0]  = A_rho[3][3][0];
   assign A_pi[3][0][1]  = A_rho[3][3][1];
   assign A_pi[3][0][2]  = A_rho[3][3][2];
   assign A_pi[3][0][3]  = A_rho[3][3][3];
   assign A_pi[3][0][4]  = A_rho[3][3][4];
   assign A_pi[3][0][5]  = A_rho[3][3][5];
   assign A_pi[3][0][6]  = A_rho[3][3][6];
   assign A_pi[3][0][7]  = A_rho[3][3][7];
   assign A_pi[3][0][8]  = A_rho[3][3][8];
   assign A_pi[3][0][9]  = A_rho[3][3][9];
   assign A_pi[3][0][10]  = A_rho[3][3][10];
   assign A_pi[3][0][11]  = A_rho[3][3][11];
   assign A_pi[3][0][12]  = A_rho[3][3][12];
   assign A_pi[3][0][13]  = A_rho[3][3][13];
   assign A_pi[3][0][14]  = A_rho[3][3][14];
   assign A_pi[3][0][15]  = A_rho[3][3][15];
   assign A_pi[3][0][16]  = A_rho[3][3][16];
   assign A_pi[3][0][17]  = A_rho[3][3][17];
   assign A_pi[3][0][18]  = A_rho[3][3][18];
   assign A_pi[3][0][19]  = A_rho[3][3][19];
   assign A_pi[3][0][20]  = A_rho[3][3][20];
   assign A_pi[3][0][21]  = A_rho[3][3][21];
   assign A_pi[3][0][22]  = A_rho[3][3][22];
   assign A_pi[3][0][23]  = A_rho[3][3][23];
   assign A_pi[3][0][24]  = A_rho[3][3][24];
   assign A_pi[3][0][25]  = A_rho[3][3][25];
   assign A_pi[3][0][26]  = A_rho[3][3][26];
   assign A_pi[3][0][27]  = A_rho[3][3][27];
   assign A_pi[3][0][28]  = A_rho[3][3][28];
   assign A_pi[3][0][29]  = A_rho[3][3][29];
   assign A_pi[3][0][30]  = A_rho[3][3][30];
   assign A_pi[3][0][31]  = A_rho[3][3][31];
   assign A_pi[3][0][32]  = A_rho[3][3][32];
   assign A_pi[3][0][33]  = A_rho[3][3][33];
   assign A_pi[3][0][34]  = A_rho[3][3][34];
   assign A_pi[3][0][35]  = A_rho[3][3][35];
   assign A_pi[3][0][36]  = A_rho[3][3][36];
   assign A_pi[3][0][37]  = A_rho[3][3][37];
   assign A_pi[3][0][38]  = A_rho[3][3][38];
   assign A_pi[3][0][39]  = A_rho[3][3][39];
   assign A_pi[3][0][40]  = A_rho[3][3][40];
   assign A_pi[3][0][41]  = A_rho[3][3][41];
   assign A_pi[3][0][42]  = A_rho[3][3][42];
   assign A_pi[3][0][43]  = A_rho[3][3][43];
   assign A_pi[3][0][44]  = A_rho[3][3][44];
   assign A_pi[3][0][45]  = A_rho[3][3][45];
   assign A_pi[3][0][46]  = A_rho[3][3][46];
   assign A_pi[3][0][47]  = A_rho[3][3][47];
   assign A_pi[3][0][48]  = A_rho[3][3][48];
   assign A_pi[3][0][49]  = A_rho[3][3][49];
   assign A_pi[3][0][50]  = A_rho[3][3][50];
   assign A_pi[3][0][51]  = A_rho[3][3][51];
   assign A_pi[3][0][52]  = A_rho[3][3][52];
   assign A_pi[3][0][53]  = A_rho[3][3][53];
   assign A_pi[3][0][54]  = A_rho[3][3][54];
   assign A_pi[3][0][55]  = A_rho[3][3][55];
   assign A_pi[3][0][56]  = A_rho[3][3][56];
   assign A_pi[3][0][57]  = A_rho[3][3][57];
   assign A_pi[3][0][58]  = A_rho[3][3][58];
   assign A_pi[3][0][59]  = A_rho[3][3][59];
   assign A_pi[3][0][60]  = A_rho[3][3][60];
   assign A_pi[3][0][61]  = A_rho[3][3][61];
   assign A_pi[3][0][62]  = A_rho[3][3][62];
   assign A_pi[3][0][63]  = A_rho[3][3][63];
   assign A_pi[3][1][0]  = A_rho[1][3][0];
   assign A_pi[3][1][1]  = A_rho[1][3][1];
   assign A_pi[3][1][2]  = A_rho[1][3][2];
   assign A_pi[3][1][3]  = A_rho[1][3][3];
   assign A_pi[3][1][4]  = A_rho[1][3][4];
   assign A_pi[3][1][5]  = A_rho[1][3][5];
   assign A_pi[3][1][6]  = A_rho[1][3][6];
   assign A_pi[3][1][7]  = A_rho[1][3][7];
   assign A_pi[3][1][8]  = A_rho[1][3][8];
   assign A_pi[3][1][9]  = A_rho[1][3][9];
   assign A_pi[3][1][10]  = A_rho[1][3][10];
   assign A_pi[3][1][11]  = A_rho[1][3][11];
   assign A_pi[3][1][12]  = A_rho[1][3][12];
   assign A_pi[3][1][13]  = A_rho[1][3][13];
   assign A_pi[3][1][14]  = A_rho[1][3][14];
   assign A_pi[3][1][15]  = A_rho[1][3][15];
   assign A_pi[3][1][16]  = A_rho[1][3][16];
   assign A_pi[3][1][17]  = A_rho[1][3][17];
   assign A_pi[3][1][18]  = A_rho[1][3][18];
   assign A_pi[3][1][19]  = A_rho[1][3][19];
   assign A_pi[3][1][20]  = A_rho[1][3][20];
   assign A_pi[3][1][21]  = A_rho[1][3][21];
   assign A_pi[3][1][22]  = A_rho[1][3][22];
   assign A_pi[3][1][23]  = A_rho[1][3][23];
   assign A_pi[3][1][24]  = A_rho[1][3][24];
   assign A_pi[3][1][25]  = A_rho[1][3][25];
   assign A_pi[3][1][26]  = A_rho[1][3][26];
   assign A_pi[3][1][27]  = A_rho[1][3][27];
   assign A_pi[3][1][28]  = A_rho[1][3][28];
   assign A_pi[3][1][29]  = A_rho[1][3][29];
   assign A_pi[3][1][30]  = A_rho[1][3][30];
   assign A_pi[3][1][31]  = A_rho[1][3][31];
   assign A_pi[3][1][32]  = A_rho[1][3][32];
   assign A_pi[3][1][33]  = A_rho[1][3][33];
   assign A_pi[3][1][34]  = A_rho[1][3][34];
   assign A_pi[3][1][35]  = A_rho[1][3][35];
   assign A_pi[3][1][36]  = A_rho[1][3][36];
   assign A_pi[3][1][37]  = A_rho[1][3][37];
   assign A_pi[3][1][38]  = A_rho[1][3][38];
   assign A_pi[3][1][39]  = A_rho[1][3][39];
   assign A_pi[3][1][40]  = A_rho[1][3][40];
   assign A_pi[3][1][41]  = A_rho[1][3][41];
   assign A_pi[3][1][42]  = A_rho[1][3][42];
   assign A_pi[3][1][43]  = A_rho[1][3][43];
   assign A_pi[3][1][44]  = A_rho[1][3][44];
   assign A_pi[3][1][45]  = A_rho[1][3][45];
   assign A_pi[3][1][46]  = A_rho[1][3][46];
   assign A_pi[3][1][47]  = A_rho[1][3][47];
   assign A_pi[3][1][48]  = A_rho[1][3][48];
   assign A_pi[3][1][49]  = A_rho[1][3][49];
   assign A_pi[3][1][50]  = A_rho[1][3][50];
   assign A_pi[3][1][51]  = A_rho[1][3][51];
   assign A_pi[3][1][52]  = A_rho[1][3][52];
   assign A_pi[3][1][53]  = A_rho[1][3][53];
   assign A_pi[3][1][54]  = A_rho[1][3][54];
   assign A_pi[3][1][55]  = A_rho[1][3][55];
   assign A_pi[3][1][56]  = A_rho[1][3][56];
   assign A_pi[3][1][57]  = A_rho[1][3][57];
   assign A_pi[3][1][58]  = A_rho[1][3][58];
   assign A_pi[3][1][59]  = A_rho[1][3][59];
   assign A_pi[3][1][60]  = A_rho[1][3][60];
   assign A_pi[3][1][61]  = A_rho[1][3][61];
   assign A_pi[3][1][62]  = A_rho[1][3][62];
   assign A_pi[3][1][63]  = A_rho[1][3][63];
   assign A_pi[3][2][0]  = A_rho[4][3][0];
   assign A_pi[3][2][1]  = A_rho[4][3][1];
   assign A_pi[3][2][2]  = A_rho[4][3][2];
   assign A_pi[3][2][3]  = A_rho[4][3][3];
   assign A_pi[3][2][4]  = A_rho[4][3][4];
   assign A_pi[3][2][5]  = A_rho[4][3][5];
   assign A_pi[3][2][6]  = A_rho[4][3][6];
   assign A_pi[3][2][7]  = A_rho[4][3][7];
   assign A_pi[3][2][8]  = A_rho[4][3][8];
   assign A_pi[3][2][9]  = A_rho[4][3][9];
   assign A_pi[3][2][10]  = A_rho[4][3][10];
   assign A_pi[3][2][11]  = A_rho[4][3][11];
   assign A_pi[3][2][12]  = A_rho[4][3][12];
   assign A_pi[3][2][13]  = A_rho[4][3][13];
   assign A_pi[3][2][14]  = A_rho[4][3][14];
   assign A_pi[3][2][15]  = A_rho[4][3][15];
   assign A_pi[3][2][16]  = A_rho[4][3][16];
   assign A_pi[3][2][17]  = A_rho[4][3][17];
   assign A_pi[3][2][18]  = A_rho[4][3][18];
   assign A_pi[3][2][19]  = A_rho[4][3][19];
   assign A_pi[3][2][20]  = A_rho[4][3][20];
   assign A_pi[3][2][21]  = A_rho[4][3][21];
   assign A_pi[3][2][22]  = A_rho[4][3][22];
   assign A_pi[3][2][23]  = A_rho[4][3][23];
   assign A_pi[3][2][24]  = A_rho[4][3][24];
   assign A_pi[3][2][25]  = A_rho[4][3][25];
   assign A_pi[3][2][26]  = A_rho[4][3][26];
   assign A_pi[3][2][27]  = A_rho[4][3][27];
   assign A_pi[3][2][28]  = A_rho[4][3][28];
   assign A_pi[3][2][29]  = A_rho[4][3][29];
   assign A_pi[3][2][30]  = A_rho[4][3][30];
   assign A_pi[3][2][31]  = A_rho[4][3][31];
   assign A_pi[3][2][32]  = A_rho[4][3][32];
   assign A_pi[3][2][33]  = A_rho[4][3][33];
   assign A_pi[3][2][34]  = A_rho[4][3][34];
   assign A_pi[3][2][35]  = A_rho[4][3][35];
   assign A_pi[3][2][36]  = A_rho[4][3][36];
   assign A_pi[3][2][37]  = A_rho[4][3][37];
   assign A_pi[3][2][38]  = A_rho[4][3][38];
   assign A_pi[3][2][39]  = A_rho[4][3][39];
   assign A_pi[3][2][40]  = A_rho[4][3][40];
   assign A_pi[3][2][41]  = A_rho[4][3][41];
   assign A_pi[3][2][42]  = A_rho[4][3][42];
   assign A_pi[3][2][43]  = A_rho[4][3][43];
   assign A_pi[3][2][44]  = A_rho[4][3][44];
   assign A_pi[3][2][45]  = A_rho[4][3][45];
   assign A_pi[3][2][46]  = A_rho[4][3][46];
   assign A_pi[3][2][47]  = A_rho[4][3][47];
   assign A_pi[3][2][48]  = A_rho[4][3][48];
   assign A_pi[3][2][49]  = A_rho[4][3][49];
   assign A_pi[3][2][50]  = A_rho[4][3][50];
   assign A_pi[3][2][51]  = A_rho[4][3][51];
   assign A_pi[3][2][52]  = A_rho[4][3][52];
   assign A_pi[3][2][53]  = A_rho[4][3][53];
   assign A_pi[3][2][54]  = A_rho[4][3][54];
   assign A_pi[3][2][55]  = A_rho[4][3][55];
   assign A_pi[3][2][56]  = A_rho[4][3][56];
   assign A_pi[3][2][57]  = A_rho[4][3][57];
   assign A_pi[3][2][58]  = A_rho[4][3][58];
   assign A_pi[3][2][59]  = A_rho[4][3][59];
   assign A_pi[3][2][60]  = A_rho[4][3][60];
   assign A_pi[3][2][61]  = A_rho[4][3][61];
   assign A_pi[3][2][62]  = A_rho[4][3][62];
   assign A_pi[3][2][63]  = A_rho[4][3][63];
   assign A_pi[3][3][0]  = A_rho[2][3][0];
   assign A_pi[3][3][1]  = A_rho[2][3][1];
   assign A_pi[3][3][2]  = A_rho[2][3][2];
   assign A_pi[3][3][3]  = A_rho[2][3][3];
   assign A_pi[3][3][4]  = A_rho[2][3][4];
   assign A_pi[3][3][5]  = A_rho[2][3][5];
   assign A_pi[3][3][6]  = A_rho[2][3][6];
   assign A_pi[3][3][7]  = A_rho[2][3][7];
   assign A_pi[3][3][8]  = A_rho[2][3][8];
   assign A_pi[3][3][9]  = A_rho[2][3][9];
   assign A_pi[3][3][10]  = A_rho[2][3][10];
   assign A_pi[3][3][11]  = A_rho[2][3][11];
   assign A_pi[3][3][12]  = A_rho[2][3][12];
   assign A_pi[3][3][13]  = A_rho[2][3][13];
   assign A_pi[3][3][14]  = A_rho[2][3][14];
   assign A_pi[3][3][15]  = A_rho[2][3][15];
   assign A_pi[3][3][16]  = A_rho[2][3][16];
   assign A_pi[3][3][17]  = A_rho[2][3][17];
   assign A_pi[3][3][18]  = A_rho[2][3][18];
   assign A_pi[3][3][19]  = A_rho[2][3][19];
   assign A_pi[3][3][20]  = A_rho[2][3][20];
   assign A_pi[3][3][21]  = A_rho[2][3][21];
   assign A_pi[3][3][22]  = A_rho[2][3][22];
   assign A_pi[3][3][23]  = A_rho[2][3][23];
   assign A_pi[3][3][24]  = A_rho[2][3][24];
   assign A_pi[3][3][25]  = A_rho[2][3][25];
   assign A_pi[3][3][26]  = A_rho[2][3][26];
   assign A_pi[3][3][27]  = A_rho[2][3][27];
   assign A_pi[3][3][28]  = A_rho[2][3][28];
   assign A_pi[3][3][29]  = A_rho[2][3][29];
   assign A_pi[3][3][30]  = A_rho[2][3][30];
   assign A_pi[3][3][31]  = A_rho[2][3][31];
   assign A_pi[3][3][32]  = A_rho[2][3][32];
   assign A_pi[3][3][33]  = A_rho[2][3][33];
   assign A_pi[3][3][34]  = A_rho[2][3][34];
   assign A_pi[3][3][35]  = A_rho[2][3][35];
   assign A_pi[3][3][36]  = A_rho[2][3][36];
   assign A_pi[3][3][37]  = A_rho[2][3][37];
   assign A_pi[3][3][38]  = A_rho[2][3][38];
   assign A_pi[3][3][39]  = A_rho[2][3][39];
   assign A_pi[3][3][40]  = A_rho[2][3][40];
   assign A_pi[3][3][41]  = A_rho[2][3][41];
   assign A_pi[3][3][42]  = A_rho[2][3][42];
   assign A_pi[3][3][43]  = A_rho[2][3][43];
   assign A_pi[3][3][44]  = A_rho[2][3][44];
   assign A_pi[3][3][45]  = A_rho[2][3][45];
   assign A_pi[3][3][46]  = A_rho[2][3][46];
   assign A_pi[3][3][47]  = A_rho[2][3][47];
   assign A_pi[3][3][48]  = A_rho[2][3][48];
   assign A_pi[3][3][49]  = A_rho[2][3][49];
   assign A_pi[3][3][50]  = A_rho[2][3][50];
   assign A_pi[3][3][51]  = A_rho[2][3][51];
   assign A_pi[3][3][52]  = A_rho[2][3][52];
   assign A_pi[3][3][53]  = A_rho[2][3][53];
   assign A_pi[3][3][54]  = A_rho[2][3][54];
   assign A_pi[3][3][55]  = A_rho[2][3][55];
   assign A_pi[3][3][56]  = A_rho[2][3][56];
   assign A_pi[3][3][57]  = A_rho[2][3][57];
   assign A_pi[3][3][58]  = A_rho[2][3][58];
   assign A_pi[3][3][59]  = A_rho[2][3][59];
   assign A_pi[3][3][60]  = A_rho[2][3][60];
   assign A_pi[3][3][61]  = A_rho[2][3][61];
   assign A_pi[3][3][62]  = A_rho[2][3][62];
   assign A_pi[3][3][63]  = A_rho[2][3][63];
   assign A_pi[3][4][0]  = A_rho[0][3][0];
   assign A_pi[3][4][1]  = A_rho[0][3][1];
   assign A_pi[3][4][2]  = A_rho[0][3][2];
   assign A_pi[3][4][3]  = A_rho[0][3][3];
   assign A_pi[3][4][4]  = A_rho[0][3][4];
   assign A_pi[3][4][5]  = A_rho[0][3][5];
   assign A_pi[3][4][6]  = A_rho[0][3][6];
   assign A_pi[3][4][7]  = A_rho[0][3][7];
   assign A_pi[3][4][8]  = A_rho[0][3][8];
   assign A_pi[3][4][9]  = A_rho[0][3][9];
   assign A_pi[3][4][10]  = A_rho[0][3][10];
   assign A_pi[3][4][11]  = A_rho[0][3][11];
   assign A_pi[3][4][12]  = A_rho[0][3][12];
   assign A_pi[3][4][13]  = A_rho[0][3][13];
   assign A_pi[3][4][14]  = A_rho[0][3][14];
   assign A_pi[3][4][15]  = A_rho[0][3][15];
   assign A_pi[3][4][16]  = A_rho[0][3][16];
   assign A_pi[3][4][17]  = A_rho[0][3][17];
   assign A_pi[3][4][18]  = A_rho[0][3][18];
   assign A_pi[3][4][19]  = A_rho[0][3][19];
   assign A_pi[3][4][20]  = A_rho[0][3][20];
   assign A_pi[3][4][21]  = A_rho[0][3][21];
   assign A_pi[3][4][22]  = A_rho[0][3][22];
   assign A_pi[3][4][23]  = A_rho[0][3][23];
   assign A_pi[3][4][24]  = A_rho[0][3][24];
   assign A_pi[3][4][25]  = A_rho[0][3][25];
   assign A_pi[3][4][26]  = A_rho[0][3][26];
   assign A_pi[3][4][27]  = A_rho[0][3][27];
   assign A_pi[3][4][28]  = A_rho[0][3][28];
   assign A_pi[3][4][29]  = A_rho[0][3][29];
   assign A_pi[3][4][30]  = A_rho[0][3][30];
   assign A_pi[3][4][31]  = A_rho[0][3][31];
   assign A_pi[3][4][32]  = A_rho[0][3][32];
   assign A_pi[3][4][33]  = A_rho[0][3][33];
   assign A_pi[3][4][34]  = A_rho[0][3][34];
   assign A_pi[3][4][35]  = A_rho[0][3][35];
   assign A_pi[3][4][36]  = A_rho[0][3][36];
   assign A_pi[3][4][37]  = A_rho[0][3][37];
   assign A_pi[3][4][38]  = A_rho[0][3][38];
   assign A_pi[3][4][39]  = A_rho[0][3][39];
   assign A_pi[3][4][40]  = A_rho[0][3][40];
   assign A_pi[3][4][41]  = A_rho[0][3][41];
   assign A_pi[3][4][42]  = A_rho[0][3][42];
   assign A_pi[3][4][43]  = A_rho[0][3][43];
   assign A_pi[3][4][44]  = A_rho[0][3][44];
   assign A_pi[3][4][45]  = A_rho[0][3][45];
   assign A_pi[3][4][46]  = A_rho[0][3][46];
   assign A_pi[3][4][47]  = A_rho[0][3][47];
   assign A_pi[3][4][48]  = A_rho[0][3][48];
   assign A_pi[3][4][49]  = A_rho[0][3][49];
   assign A_pi[3][4][50]  = A_rho[0][3][50];
   assign A_pi[3][4][51]  = A_rho[0][3][51];
   assign A_pi[3][4][52]  = A_rho[0][3][52];
   assign A_pi[3][4][53]  = A_rho[0][3][53];
   assign A_pi[3][4][54]  = A_rho[0][3][54];
   assign A_pi[3][4][55]  = A_rho[0][3][55];
   assign A_pi[3][4][56]  = A_rho[0][3][56];
   assign A_pi[3][4][57]  = A_rho[0][3][57];
   assign A_pi[3][4][58]  = A_rho[0][3][58];
   assign A_pi[3][4][59]  = A_rho[0][3][59];
   assign A_pi[3][4][60]  = A_rho[0][3][60];
   assign A_pi[3][4][61]  = A_rho[0][3][61];
   assign A_pi[3][4][62]  = A_rho[0][3][62];
   assign A_pi[3][4][63]  = A_rho[0][3][63];
   assign A_pi[4][0][0]  = A_rho[4][4][0];
   assign A_pi[4][0][1]  = A_rho[4][4][1];
   assign A_pi[4][0][2]  = A_rho[4][4][2];
   assign A_pi[4][0][3]  = A_rho[4][4][3];
   assign A_pi[4][0][4]  = A_rho[4][4][4];
   assign A_pi[4][0][5]  = A_rho[4][4][5];
   assign A_pi[4][0][6]  = A_rho[4][4][6];
   assign A_pi[4][0][7]  = A_rho[4][4][7];
   assign A_pi[4][0][8]  = A_rho[4][4][8];
   assign A_pi[4][0][9]  = A_rho[4][4][9];
   assign A_pi[4][0][10]  = A_rho[4][4][10];
   assign A_pi[4][0][11]  = A_rho[4][4][11];
   assign A_pi[4][0][12]  = A_rho[4][4][12];
   assign A_pi[4][0][13]  = A_rho[4][4][13];
   assign A_pi[4][0][14]  = A_rho[4][4][14];
   assign A_pi[4][0][15]  = A_rho[4][4][15];
   assign A_pi[4][0][16]  = A_rho[4][4][16];
   assign A_pi[4][0][17]  = A_rho[4][4][17];
   assign A_pi[4][0][18]  = A_rho[4][4][18];
   assign A_pi[4][0][19]  = A_rho[4][4][19];
   assign A_pi[4][0][20]  = A_rho[4][4][20];
   assign A_pi[4][0][21]  = A_rho[4][4][21];
   assign A_pi[4][0][22]  = A_rho[4][4][22];
   assign A_pi[4][0][23]  = A_rho[4][4][23];
   assign A_pi[4][0][24]  = A_rho[4][4][24];
   assign A_pi[4][0][25]  = A_rho[4][4][25];
   assign A_pi[4][0][26]  = A_rho[4][4][26];
   assign A_pi[4][0][27]  = A_rho[4][4][27];
   assign A_pi[4][0][28]  = A_rho[4][4][28];
   assign A_pi[4][0][29]  = A_rho[4][4][29];
   assign A_pi[4][0][30]  = A_rho[4][4][30];
   assign A_pi[4][0][31]  = A_rho[4][4][31];
   assign A_pi[4][0][32]  = A_rho[4][4][32];
   assign A_pi[4][0][33]  = A_rho[4][4][33];
   assign A_pi[4][0][34]  = A_rho[4][4][34];
   assign A_pi[4][0][35]  = A_rho[4][4][35];
   assign A_pi[4][0][36]  = A_rho[4][4][36];
   assign A_pi[4][0][37]  = A_rho[4][4][37];
   assign A_pi[4][0][38]  = A_rho[4][4][38];
   assign A_pi[4][0][39]  = A_rho[4][4][39];
   assign A_pi[4][0][40]  = A_rho[4][4][40];
   assign A_pi[4][0][41]  = A_rho[4][4][41];
   assign A_pi[4][0][42]  = A_rho[4][4][42];
   assign A_pi[4][0][43]  = A_rho[4][4][43];
   assign A_pi[4][0][44]  = A_rho[4][4][44];
   assign A_pi[4][0][45]  = A_rho[4][4][45];
   assign A_pi[4][0][46]  = A_rho[4][4][46];
   assign A_pi[4][0][47]  = A_rho[4][4][47];
   assign A_pi[4][0][48]  = A_rho[4][4][48];
   assign A_pi[4][0][49]  = A_rho[4][4][49];
   assign A_pi[4][0][50]  = A_rho[4][4][50];
   assign A_pi[4][0][51]  = A_rho[4][4][51];
   assign A_pi[4][0][52]  = A_rho[4][4][52];
   assign A_pi[4][0][53]  = A_rho[4][4][53];
   assign A_pi[4][0][54]  = A_rho[4][4][54];
   assign A_pi[4][0][55]  = A_rho[4][4][55];
   assign A_pi[4][0][56]  = A_rho[4][4][56];
   assign A_pi[4][0][57]  = A_rho[4][4][57];
   assign A_pi[4][0][58]  = A_rho[4][4][58];
   assign A_pi[4][0][59]  = A_rho[4][4][59];
   assign A_pi[4][0][60]  = A_rho[4][4][60];
   assign A_pi[4][0][61]  = A_rho[4][4][61];
   assign A_pi[4][0][62]  = A_rho[4][4][62];
   assign A_pi[4][0][63]  = A_rho[4][4][63];
   assign A_pi[4][1][0]  = A_rho[2][4][0];
   assign A_pi[4][1][1]  = A_rho[2][4][1];
   assign A_pi[4][1][2]  = A_rho[2][4][2];
   assign A_pi[4][1][3]  = A_rho[2][4][3];
   assign A_pi[4][1][4]  = A_rho[2][4][4];
   assign A_pi[4][1][5]  = A_rho[2][4][5];
   assign A_pi[4][1][6]  = A_rho[2][4][6];
   assign A_pi[4][1][7]  = A_rho[2][4][7];
   assign A_pi[4][1][8]  = A_rho[2][4][8];
   assign A_pi[4][1][9]  = A_rho[2][4][9];
   assign A_pi[4][1][10]  = A_rho[2][4][10];
   assign A_pi[4][1][11]  = A_rho[2][4][11];
   assign A_pi[4][1][12]  = A_rho[2][4][12];
   assign A_pi[4][1][13]  = A_rho[2][4][13];
   assign A_pi[4][1][14]  = A_rho[2][4][14];
   assign A_pi[4][1][15]  = A_rho[2][4][15];
   assign A_pi[4][1][16]  = A_rho[2][4][16];
   assign A_pi[4][1][17]  = A_rho[2][4][17];
   assign A_pi[4][1][18]  = A_rho[2][4][18];
   assign A_pi[4][1][19]  = A_rho[2][4][19];
   assign A_pi[4][1][20]  = A_rho[2][4][20];
   assign A_pi[4][1][21]  = A_rho[2][4][21];
   assign A_pi[4][1][22]  = A_rho[2][4][22];
   assign A_pi[4][1][23]  = A_rho[2][4][23];
   assign A_pi[4][1][24]  = A_rho[2][4][24];
   assign A_pi[4][1][25]  = A_rho[2][4][25];
   assign A_pi[4][1][26]  = A_rho[2][4][26];
   assign A_pi[4][1][27]  = A_rho[2][4][27];
   assign A_pi[4][1][28]  = A_rho[2][4][28];
   assign A_pi[4][1][29]  = A_rho[2][4][29];
   assign A_pi[4][1][30]  = A_rho[2][4][30];
   assign A_pi[4][1][31]  = A_rho[2][4][31];
   assign A_pi[4][1][32]  = A_rho[2][4][32];
   assign A_pi[4][1][33]  = A_rho[2][4][33];
   assign A_pi[4][1][34]  = A_rho[2][4][34];
   assign A_pi[4][1][35]  = A_rho[2][4][35];
   assign A_pi[4][1][36]  = A_rho[2][4][36];
   assign A_pi[4][1][37]  = A_rho[2][4][37];
   assign A_pi[4][1][38]  = A_rho[2][4][38];
   assign A_pi[4][1][39]  = A_rho[2][4][39];
   assign A_pi[4][1][40]  = A_rho[2][4][40];
   assign A_pi[4][1][41]  = A_rho[2][4][41];
   assign A_pi[4][1][42]  = A_rho[2][4][42];
   assign A_pi[4][1][43]  = A_rho[2][4][43];
   assign A_pi[4][1][44]  = A_rho[2][4][44];
   assign A_pi[4][1][45]  = A_rho[2][4][45];
   assign A_pi[4][1][46]  = A_rho[2][4][46];
   assign A_pi[4][1][47]  = A_rho[2][4][47];
   assign A_pi[4][1][48]  = A_rho[2][4][48];
   assign A_pi[4][1][49]  = A_rho[2][4][49];
   assign A_pi[4][1][50]  = A_rho[2][4][50];
   assign A_pi[4][1][51]  = A_rho[2][4][51];
   assign A_pi[4][1][52]  = A_rho[2][4][52];
   assign A_pi[4][1][53]  = A_rho[2][4][53];
   assign A_pi[4][1][54]  = A_rho[2][4][54];
   assign A_pi[4][1][55]  = A_rho[2][4][55];
   assign A_pi[4][1][56]  = A_rho[2][4][56];
   assign A_pi[4][1][57]  = A_rho[2][4][57];
   assign A_pi[4][1][58]  = A_rho[2][4][58];
   assign A_pi[4][1][59]  = A_rho[2][4][59];
   assign A_pi[4][1][60]  = A_rho[2][4][60];
   assign A_pi[4][1][61]  = A_rho[2][4][61];
   assign A_pi[4][1][62]  = A_rho[2][4][62];
   assign A_pi[4][1][63]  = A_rho[2][4][63];
   assign A_pi[4][2][0]  = A_rho[0][4][0];
   assign A_pi[4][2][1]  = A_rho[0][4][1];
   assign A_pi[4][2][2]  = A_rho[0][4][2];
   assign A_pi[4][2][3]  = A_rho[0][4][3];
   assign A_pi[4][2][4]  = A_rho[0][4][4];
   assign A_pi[4][2][5]  = A_rho[0][4][5];
   assign A_pi[4][2][6]  = A_rho[0][4][6];
   assign A_pi[4][2][7]  = A_rho[0][4][7];
   assign A_pi[4][2][8]  = A_rho[0][4][8];
   assign A_pi[4][2][9]  = A_rho[0][4][9];
   assign A_pi[4][2][10]  = A_rho[0][4][10];
   assign A_pi[4][2][11]  = A_rho[0][4][11];
   assign A_pi[4][2][12]  = A_rho[0][4][12];
   assign A_pi[4][2][13]  = A_rho[0][4][13];
   assign A_pi[4][2][14]  = A_rho[0][4][14];
   assign A_pi[4][2][15]  = A_rho[0][4][15];
   assign A_pi[4][2][16]  = A_rho[0][4][16];
   assign A_pi[4][2][17]  = A_rho[0][4][17];
   assign A_pi[4][2][18]  = A_rho[0][4][18];
   assign A_pi[4][2][19]  = A_rho[0][4][19];
   assign A_pi[4][2][20]  = A_rho[0][4][20];
   assign A_pi[4][2][21]  = A_rho[0][4][21];
   assign A_pi[4][2][22]  = A_rho[0][4][22];
   assign A_pi[4][2][23]  = A_rho[0][4][23];
   assign A_pi[4][2][24]  = A_rho[0][4][24];
   assign A_pi[4][2][25]  = A_rho[0][4][25];
   assign A_pi[4][2][26]  = A_rho[0][4][26];
   assign A_pi[4][2][27]  = A_rho[0][4][27];
   assign A_pi[4][2][28]  = A_rho[0][4][28];
   assign A_pi[4][2][29]  = A_rho[0][4][29];
   assign A_pi[4][2][30]  = A_rho[0][4][30];
   assign A_pi[4][2][31]  = A_rho[0][4][31];
   assign A_pi[4][2][32]  = A_rho[0][4][32];
   assign A_pi[4][2][33]  = A_rho[0][4][33];
   assign A_pi[4][2][34]  = A_rho[0][4][34];
   assign A_pi[4][2][35]  = A_rho[0][4][35];
   assign A_pi[4][2][36]  = A_rho[0][4][36];
   assign A_pi[4][2][37]  = A_rho[0][4][37];
   assign A_pi[4][2][38]  = A_rho[0][4][38];
   assign A_pi[4][2][39]  = A_rho[0][4][39];
   assign A_pi[4][2][40]  = A_rho[0][4][40];
   assign A_pi[4][2][41]  = A_rho[0][4][41];
   assign A_pi[4][2][42]  = A_rho[0][4][42];
   assign A_pi[4][2][43]  = A_rho[0][4][43];
   assign A_pi[4][2][44]  = A_rho[0][4][44];
   assign A_pi[4][2][45]  = A_rho[0][4][45];
   assign A_pi[4][2][46]  = A_rho[0][4][46];
   assign A_pi[4][2][47]  = A_rho[0][4][47];
   assign A_pi[4][2][48]  = A_rho[0][4][48];
   assign A_pi[4][2][49]  = A_rho[0][4][49];
   assign A_pi[4][2][50]  = A_rho[0][4][50];
   assign A_pi[4][2][51]  = A_rho[0][4][51];
   assign A_pi[4][2][52]  = A_rho[0][4][52];
   assign A_pi[4][2][53]  = A_rho[0][4][53];
   assign A_pi[4][2][54]  = A_rho[0][4][54];
   assign A_pi[4][2][55]  = A_rho[0][4][55];
   assign A_pi[4][2][56]  = A_rho[0][4][56];
   assign A_pi[4][2][57]  = A_rho[0][4][57];
   assign A_pi[4][2][58]  = A_rho[0][4][58];
   assign A_pi[4][2][59]  = A_rho[0][4][59];
   assign A_pi[4][2][60]  = A_rho[0][4][60];
   assign A_pi[4][2][61]  = A_rho[0][4][61];
   assign A_pi[4][2][62]  = A_rho[0][4][62];
   assign A_pi[4][2][63]  = A_rho[0][4][63];
   assign A_pi[4][3][0]  = A_rho[3][4][0];
   assign A_pi[4][3][1]  = A_rho[3][4][1];
   assign A_pi[4][3][2]  = A_rho[3][4][2];
   assign A_pi[4][3][3]  = A_rho[3][4][3];
   assign A_pi[4][3][4]  = A_rho[3][4][4];
   assign A_pi[4][3][5]  = A_rho[3][4][5];
   assign A_pi[4][3][6]  = A_rho[3][4][6];
   assign A_pi[4][3][7]  = A_rho[3][4][7];
   assign A_pi[4][3][8]  = A_rho[3][4][8];
   assign A_pi[4][3][9]  = A_rho[3][4][9];
   assign A_pi[4][3][10]  = A_rho[3][4][10];
   assign A_pi[4][3][11]  = A_rho[3][4][11];
   assign A_pi[4][3][12]  = A_rho[3][4][12];
   assign A_pi[4][3][13]  = A_rho[3][4][13];
   assign A_pi[4][3][14]  = A_rho[3][4][14];
   assign A_pi[4][3][15]  = A_rho[3][4][15];
   assign A_pi[4][3][16]  = A_rho[3][4][16];
   assign A_pi[4][3][17]  = A_rho[3][4][17];
   assign A_pi[4][3][18]  = A_rho[3][4][18];
   assign A_pi[4][3][19]  = A_rho[3][4][19];
   assign A_pi[4][3][20]  = A_rho[3][4][20];
   assign A_pi[4][3][21]  = A_rho[3][4][21];
   assign A_pi[4][3][22]  = A_rho[3][4][22];
   assign A_pi[4][3][23]  = A_rho[3][4][23];
   assign A_pi[4][3][24]  = A_rho[3][4][24];
   assign A_pi[4][3][25]  = A_rho[3][4][25];
   assign A_pi[4][3][26]  = A_rho[3][4][26];
   assign A_pi[4][3][27]  = A_rho[3][4][27];
   assign A_pi[4][3][28]  = A_rho[3][4][28];
   assign A_pi[4][3][29]  = A_rho[3][4][29];
   assign A_pi[4][3][30]  = A_rho[3][4][30];
   assign A_pi[4][3][31]  = A_rho[3][4][31];
   assign A_pi[4][3][32]  = A_rho[3][4][32];
   assign A_pi[4][3][33]  = A_rho[3][4][33];
   assign A_pi[4][3][34]  = A_rho[3][4][34];
   assign A_pi[4][3][35]  = A_rho[3][4][35];
   assign A_pi[4][3][36]  = A_rho[3][4][36];
   assign A_pi[4][3][37]  = A_rho[3][4][37];
   assign A_pi[4][3][38]  = A_rho[3][4][38];
   assign A_pi[4][3][39]  = A_rho[3][4][39];
   assign A_pi[4][3][40]  = A_rho[3][4][40];
   assign A_pi[4][3][41]  = A_rho[3][4][41];
   assign A_pi[4][3][42]  = A_rho[3][4][42];
   assign A_pi[4][3][43]  = A_rho[3][4][43];
   assign A_pi[4][3][44]  = A_rho[3][4][44];
   assign A_pi[4][3][45]  = A_rho[3][4][45];
   assign A_pi[4][3][46]  = A_rho[3][4][46];
   assign A_pi[4][3][47]  = A_rho[3][4][47];
   assign A_pi[4][3][48]  = A_rho[3][4][48];
   assign A_pi[4][3][49]  = A_rho[3][4][49];
   assign A_pi[4][3][50]  = A_rho[3][4][50];
   assign A_pi[4][3][51]  = A_rho[3][4][51];
   assign A_pi[4][3][52]  = A_rho[3][4][52];
   assign A_pi[4][3][53]  = A_rho[3][4][53];
   assign A_pi[4][3][54]  = A_rho[3][4][54];
   assign A_pi[4][3][55]  = A_rho[3][4][55];
   assign A_pi[4][3][56]  = A_rho[3][4][56];
   assign A_pi[4][3][57]  = A_rho[3][4][57];
   assign A_pi[4][3][58]  = A_rho[3][4][58];
   assign A_pi[4][3][59]  = A_rho[3][4][59];
   assign A_pi[4][3][60]  = A_rho[3][4][60];
   assign A_pi[4][3][61]  = A_rho[3][4][61];
   assign A_pi[4][3][62]  = A_rho[3][4][62];
   assign A_pi[4][3][63]  = A_rho[3][4][63];
   assign A_pi[4][4][0]  = A_rho[1][4][0];
   assign A_pi[4][4][1]  = A_rho[1][4][1];
   assign A_pi[4][4][2]  = A_rho[1][4][2];
   assign A_pi[4][4][3]  = A_rho[1][4][3];
   assign A_pi[4][4][4]  = A_rho[1][4][4];
   assign A_pi[4][4][5]  = A_rho[1][4][5];
   assign A_pi[4][4][6]  = A_rho[1][4][6];
   assign A_pi[4][4][7]  = A_rho[1][4][7];
   assign A_pi[4][4][8]  = A_rho[1][4][8];
   assign A_pi[4][4][9]  = A_rho[1][4][9];
   assign A_pi[4][4][10]  = A_rho[1][4][10];
   assign A_pi[4][4][11]  = A_rho[1][4][11];
   assign A_pi[4][4][12]  = A_rho[1][4][12];
   assign A_pi[4][4][13]  = A_rho[1][4][13];
   assign A_pi[4][4][14]  = A_rho[1][4][14];
   assign A_pi[4][4][15]  = A_rho[1][4][15];
   assign A_pi[4][4][16]  = A_rho[1][4][16];
   assign A_pi[4][4][17]  = A_rho[1][4][17];
   assign A_pi[4][4][18]  = A_rho[1][4][18];
   assign A_pi[4][4][19]  = A_rho[1][4][19];
   assign A_pi[4][4][20]  = A_rho[1][4][20];
   assign A_pi[4][4][21]  = A_rho[1][4][21];
   assign A_pi[4][4][22]  = A_rho[1][4][22];
   assign A_pi[4][4][23]  = A_rho[1][4][23];
   assign A_pi[4][4][24]  = A_rho[1][4][24];
   assign A_pi[4][4][25]  = A_rho[1][4][25];
   assign A_pi[4][4][26]  = A_rho[1][4][26];
   assign A_pi[4][4][27]  = A_rho[1][4][27];
   assign A_pi[4][4][28]  = A_rho[1][4][28];
   assign A_pi[4][4][29]  = A_rho[1][4][29];
   assign A_pi[4][4][30]  = A_rho[1][4][30];
   assign A_pi[4][4][31]  = A_rho[1][4][31];
   assign A_pi[4][4][32]  = A_rho[1][4][32];
   assign A_pi[4][4][33]  = A_rho[1][4][33];
   assign A_pi[4][4][34]  = A_rho[1][4][34];
   assign A_pi[4][4][35]  = A_rho[1][4][35];
   assign A_pi[4][4][36]  = A_rho[1][4][36];
   assign A_pi[4][4][37]  = A_rho[1][4][37];
   assign A_pi[4][4][38]  = A_rho[1][4][38];
   assign A_pi[4][4][39]  = A_rho[1][4][39];
   assign A_pi[4][4][40]  = A_rho[1][4][40];
   assign A_pi[4][4][41]  = A_rho[1][4][41];
   assign A_pi[4][4][42]  = A_rho[1][4][42];
   assign A_pi[4][4][43]  = A_rho[1][4][43];
   assign A_pi[4][4][44]  = A_rho[1][4][44];
   assign A_pi[4][4][45]  = A_rho[1][4][45];
   assign A_pi[4][4][46]  = A_rho[1][4][46];
   assign A_pi[4][4][47]  = A_rho[1][4][47];
   assign A_pi[4][4][48]  = A_rho[1][4][48];
   assign A_pi[4][4][49]  = A_rho[1][4][49];
   assign A_pi[4][4][50]  = A_rho[1][4][50];
   assign A_pi[4][4][51]  = A_rho[1][4][51];
   assign A_pi[4][4][52]  = A_rho[1][4][52];
   assign A_pi[4][4][53]  = A_rho[1][4][53];
   assign A_pi[4][4][54]  = A_rho[1][4][54];
   assign A_pi[4][4][55]  = A_rho[1][4][55];
   assign A_pi[4][4][56]  = A_rho[1][4][56];
   assign A_pi[4][4][57]  = A_rho[1][4][57];
   assign A_pi[4][4][58]  = A_rho[1][4][58];
   assign A_pi[4][4][59]  = A_rho[1][4][59];
   assign A_pi[4][4][60]  = A_rho[1][4][60];
   assign A_pi[4][4][61]  = A_rho[1][4][61];
   assign A_pi[4][4][62]  = A_rho[1][4][62];
   assign A_pi[4][4][63]  = A_rho[1][4][63];
//--------------------------- CHI ---------------------------
   assign A_chi[0][0][0]     = A[0][0][0] ^ ((~A[1][0][0]) & A[2][0][0]);
   assign A_chi[0][0][1]     = A[0][0][1] ^ ((~A[1][0][1]) & A[2][0][1]);
   assign A_chi[0][0][2]     = A[0][0][2] ^ ((~A[1][0][2]) & A[2][0][2]);
   assign A_chi[0][0][3]     = A[0][0][3] ^ ((~A[1][0][3]) & A[2][0][3]);
   assign A_chi[0][0][4]     = A[0][0][4] ^ ((~A[1][0][4]) & A[2][0][4]);
   assign A_chi[0][0][5]     = A[0][0][5] ^ ((~A[1][0][5]) & A[2][0][5]);
   assign A_chi[0][0][6]     = A[0][0][6] ^ ((~A[1][0][6]) & A[2][0][6]);
   assign A_chi[0][0][7]     = A[0][0][7] ^ ((~A[1][0][7]) & A[2][0][7]);
   assign A_chi[0][0][8]     = A[0][0][8] ^ ((~A[1][0][8]) & A[2][0][8]);
   assign A_chi[0][0][9]     = A[0][0][9] ^ ((~A[1][0][9]) & A[2][0][9]);
   assign A_chi[0][0][10]     = A[0][0][10] ^ ((~A[1][0][10]) & A[2][0][10]);
   assign A_chi[0][0][11]     = A[0][0][11] ^ ((~A[1][0][11]) & A[2][0][11]);
   assign A_chi[0][0][12]     = A[0][0][12] ^ ((~A[1][0][12]) & A[2][0][12]);
   assign A_chi[0][0][13]     = A[0][0][13] ^ ((~A[1][0][13]) & A[2][0][13]);
   assign A_chi[0][0][14]     = A[0][0][14] ^ ((~A[1][0][14]) & A[2][0][14]);
   assign A_chi[0][0][15]     = A[0][0][15] ^ ((~A[1][0][15]) & A[2][0][15]);
   assign A_chi[0][0][16]     = A[0][0][16] ^ ((~A[1][0][16]) & A[2][0][16]);
   assign A_chi[0][0][17]     = A[0][0][17] ^ ((~A[1][0][17]) & A[2][0][17]);
   assign A_chi[0][0][18]     = A[0][0][18] ^ ((~A[1][0][18]) & A[2][0][18]);
   assign A_chi[0][0][19]     = A[0][0][19] ^ ((~A[1][0][19]) & A[2][0][19]);
   assign A_chi[0][0][20]     = A[0][0][20] ^ ((~A[1][0][20]) & A[2][0][20]);
   assign A_chi[0][0][21]     = A[0][0][21] ^ ((~A[1][0][21]) & A[2][0][21]);
   assign A_chi[0][0][22]     = A[0][0][22] ^ ((~A[1][0][22]) & A[2][0][22]);
   assign A_chi[0][0][23]     = A[0][0][23] ^ ((~A[1][0][23]) & A[2][0][23]);
   assign A_chi[0][0][24]     = A[0][0][24] ^ ((~A[1][0][24]) & A[2][0][24]);
   assign A_chi[0][0][25]     = A[0][0][25] ^ ((~A[1][0][25]) & A[2][0][25]);
   assign A_chi[0][0][26]     = A[0][0][26] ^ ((~A[1][0][26]) & A[2][0][26]);
   assign A_chi[0][0][27]     = A[0][0][27] ^ ((~A[1][0][27]) & A[2][0][27]);
   assign A_chi[0][0][28]     = A[0][0][28] ^ ((~A[1][0][28]) & A[2][0][28]);
   assign A_chi[0][0][29]     = A[0][0][29] ^ ((~A[1][0][29]) & A[2][0][29]);
   assign A_chi[0][0][30]     = A[0][0][30] ^ ((~A[1][0][30]) & A[2][0][30]);
   assign A_chi[0][0][31]     = A[0][0][31] ^ ((~A[1][0][31]) & A[2][0][31]);
   assign A_chi[0][0][32]     = A[0][0][32] ^ ((~A[1][0][32]) & A[2][0][32]);
   assign A_chi[0][0][33]     = A[0][0][33] ^ ((~A[1][0][33]) & A[2][0][33]);
   assign A_chi[0][0][34]     = A[0][0][34] ^ ((~A[1][0][34]) & A[2][0][34]);
   assign A_chi[0][0][35]     = A[0][0][35] ^ ((~A[1][0][35]) & A[2][0][35]);
   assign A_chi[0][0][36]     = A[0][0][36] ^ ((~A[1][0][36]) & A[2][0][36]);
   assign A_chi[0][0][37]     = A[0][0][37] ^ ((~A[1][0][37]) & A[2][0][37]);
   assign A_chi[0][0][38]     = A[0][0][38] ^ ((~A[1][0][38]) & A[2][0][38]);
   assign A_chi[0][0][39]     = A[0][0][39] ^ ((~A[1][0][39]) & A[2][0][39]);
   assign A_chi[0][0][40]     = A[0][0][40] ^ ((~A[1][0][40]) & A[2][0][40]);
   assign A_chi[0][0][41]     = A[0][0][41] ^ ((~A[1][0][41]) & A[2][0][41]);
   assign A_chi[0][0][42]     = A[0][0][42] ^ ((~A[1][0][42]) & A[2][0][42]);
   assign A_chi[0][0][43]     = A[0][0][43] ^ ((~A[1][0][43]) & A[2][0][43]);
   assign A_chi[0][0][44]     = A[0][0][44] ^ ((~A[1][0][44]) & A[2][0][44]);
   assign A_chi[0][0][45]     = A[0][0][45] ^ ((~A[1][0][45]) & A[2][0][45]);
   assign A_chi[0][0][46]     = A[0][0][46] ^ ((~A[1][0][46]) & A[2][0][46]);
   assign A_chi[0][0][47]     = A[0][0][47] ^ ((~A[1][0][47]) & A[2][0][47]);
   assign A_chi[0][0][48]     = A[0][0][48] ^ ((~A[1][0][48]) & A[2][0][48]);
   assign A_chi[0][0][49]     = A[0][0][49] ^ ((~A[1][0][49]) & A[2][0][49]);
   assign A_chi[0][0][50]     = A[0][0][50] ^ ((~A[1][0][50]) & A[2][0][50]);
   assign A_chi[0][0][51]     = A[0][0][51] ^ ((~A[1][0][51]) & A[2][0][51]);
   assign A_chi[0][0][52]     = A[0][0][52] ^ ((~A[1][0][52]) & A[2][0][52]);
   assign A_chi[0][0][53]     = A[0][0][53] ^ ((~A[1][0][53]) & A[2][0][53]);
   assign A_chi[0][0][54]     = A[0][0][54] ^ ((~A[1][0][54]) & A[2][0][54]);
   assign A_chi[0][0][55]     = A[0][0][55] ^ ((~A[1][0][55]) & A[2][0][55]);
   assign A_chi[0][0][56]     = A[0][0][56] ^ ((~A[1][0][56]) & A[2][0][56]);
   assign A_chi[0][0][57]     = A[0][0][57] ^ ((~A[1][0][57]) & A[2][0][57]);
   assign A_chi[0][0][58]     = A[0][0][58] ^ ((~A[1][0][58]) & A[2][0][58]);
   assign A_chi[0][0][59]     = A[0][0][59] ^ ((~A[1][0][59]) & A[2][0][59]);
   assign A_chi[0][0][60]     = A[0][0][60] ^ ((~A[1][0][60]) & A[2][0][60]);
   assign A_chi[0][0][61]     = A[0][0][61] ^ ((~A[1][0][61]) & A[2][0][61]);
   assign A_chi[0][0][62]     = A[0][0][62] ^ ((~A[1][0][62]) & A[2][0][62]);
   assign A_chi[0][0][63]     = A[0][0][63] ^ ((~A[1][0][63]) & A[2][0][63]);
   assign A_chi[0][1][0]     = A[1][0][0] ^ ((~A[2][0][0]) & A[3][0][0]);
   assign A_chi[0][1][1]     = A[1][0][1] ^ ((~A[2][0][1]) & A[3][0][1]);
   assign A_chi[0][1][2]     = A[1][0][2] ^ ((~A[2][0][2]) & A[3][0][2]);
   assign A_chi[0][1][3]     = A[1][0][3] ^ ((~A[2][0][3]) & A[3][0][3]);
   assign A_chi[0][1][4]     = A[1][0][4] ^ ((~A[2][0][4]) & A[3][0][4]);
   assign A_chi[0][1][5]     = A[1][0][5] ^ ((~A[2][0][5]) & A[3][0][5]);
   assign A_chi[0][1][6]     = A[1][0][6] ^ ((~A[2][0][6]) & A[3][0][6]);
   assign A_chi[0][1][7]     = A[1][0][7] ^ ((~A[2][0][7]) & A[3][0][7]);
   assign A_chi[0][1][8]     = A[1][0][8] ^ ((~A[2][0][8]) & A[3][0][8]);
   assign A_chi[0][1][9]     = A[1][0][9] ^ ((~A[2][0][9]) & A[3][0][9]);
   assign A_chi[0][1][10]     = A[1][0][10] ^ ((~A[2][0][10]) & A[3][0][10]);
   assign A_chi[0][1][11]     = A[1][0][11] ^ ((~A[2][0][11]) & A[3][0][11]);
   assign A_chi[0][1][12]     = A[1][0][12] ^ ((~A[2][0][12]) & A[3][0][12]);
   assign A_chi[0][1][13]     = A[1][0][13] ^ ((~A[2][0][13]) & A[3][0][13]);
   assign A_chi[0][1][14]     = A[1][0][14] ^ ((~A[2][0][14]) & A[3][0][14]);
   assign A_chi[0][1][15]     = A[1][0][15] ^ ((~A[2][0][15]) & A[3][0][15]);
   assign A_chi[0][1][16]     = A[1][0][16] ^ ((~A[2][0][16]) & A[3][0][16]);
   assign A_chi[0][1][17]     = A[1][0][17] ^ ((~A[2][0][17]) & A[3][0][17]);
   assign A_chi[0][1][18]     = A[1][0][18] ^ ((~A[2][0][18]) & A[3][0][18]);
   assign A_chi[0][1][19]     = A[1][0][19] ^ ((~A[2][0][19]) & A[3][0][19]);
   assign A_chi[0][1][20]     = A[1][0][20] ^ ((~A[2][0][20]) & A[3][0][20]);
   assign A_chi[0][1][21]     = A[1][0][21] ^ ((~A[2][0][21]) & A[3][0][21]);
   assign A_chi[0][1][22]     = A[1][0][22] ^ ((~A[2][0][22]) & A[3][0][22]);
   assign A_chi[0][1][23]     = A[1][0][23] ^ ((~A[2][0][23]) & A[3][0][23]);
   assign A_chi[0][1][24]     = A[1][0][24] ^ ((~A[2][0][24]) & A[3][0][24]);
   assign A_chi[0][1][25]     = A[1][0][25] ^ ((~A[2][0][25]) & A[3][0][25]);
   assign A_chi[0][1][26]     = A[1][0][26] ^ ((~A[2][0][26]) & A[3][0][26]);
   assign A_chi[0][1][27]     = A[1][0][27] ^ ((~A[2][0][27]) & A[3][0][27]);
   assign A_chi[0][1][28]     = A[1][0][28] ^ ((~A[2][0][28]) & A[3][0][28]);
   assign A_chi[0][1][29]     = A[1][0][29] ^ ((~A[2][0][29]) & A[3][0][29]);
   assign A_chi[0][1][30]     = A[1][0][30] ^ ((~A[2][0][30]) & A[3][0][30]);
   assign A_chi[0][1][31]     = A[1][0][31] ^ ((~A[2][0][31]) & A[3][0][31]);
   assign A_chi[0][1][32]     = A[1][0][32] ^ ((~A[2][0][32]) & A[3][0][32]);
   assign A_chi[0][1][33]     = A[1][0][33] ^ ((~A[2][0][33]) & A[3][0][33]);
   assign A_chi[0][1][34]     = A[1][0][34] ^ ((~A[2][0][34]) & A[3][0][34]);
   assign A_chi[0][1][35]     = A[1][0][35] ^ ((~A[2][0][35]) & A[3][0][35]);
   assign A_chi[0][1][36]     = A[1][0][36] ^ ((~A[2][0][36]) & A[3][0][36]);
   assign A_chi[0][1][37]     = A[1][0][37] ^ ((~A[2][0][37]) & A[3][0][37]);
   assign A_chi[0][1][38]     = A[1][0][38] ^ ((~A[2][0][38]) & A[3][0][38]);
   assign A_chi[0][1][39]     = A[1][0][39] ^ ((~A[2][0][39]) & A[3][0][39]);
   assign A_chi[0][1][40]     = A[1][0][40] ^ ((~A[2][0][40]) & A[3][0][40]);
   assign A_chi[0][1][41]     = A[1][0][41] ^ ((~A[2][0][41]) & A[3][0][41]);
   assign A_chi[0][1][42]     = A[1][0][42] ^ ((~A[2][0][42]) & A[3][0][42]);
   assign A_chi[0][1][43]     = A[1][0][43] ^ ((~A[2][0][43]) & A[3][0][43]);
   assign A_chi[0][1][44]     = A[1][0][44] ^ ((~A[2][0][44]) & A[3][0][44]);
   assign A_chi[0][1][45]     = A[1][0][45] ^ ((~A[2][0][45]) & A[3][0][45]);
   assign A_chi[0][1][46]     = A[1][0][46] ^ ((~A[2][0][46]) & A[3][0][46]);
   assign A_chi[0][1][47]     = A[1][0][47] ^ ((~A[2][0][47]) & A[3][0][47]);
   assign A_chi[0][1][48]     = A[1][0][48] ^ ((~A[2][0][48]) & A[3][0][48]);
   assign A_chi[0][1][49]     = A[1][0][49] ^ ((~A[2][0][49]) & A[3][0][49]);
   assign A_chi[0][1][50]     = A[1][0][50] ^ ((~A[2][0][50]) & A[3][0][50]);
   assign A_chi[0][1][51]     = A[1][0][51] ^ ((~A[2][0][51]) & A[3][0][51]);
   assign A_chi[0][1][52]     = A[1][0][52] ^ ((~A[2][0][52]) & A[3][0][52]);
   assign A_chi[0][1][53]     = A[1][0][53] ^ ((~A[2][0][53]) & A[3][0][53]);
   assign A_chi[0][1][54]     = A[1][0][54] ^ ((~A[2][0][54]) & A[3][0][54]);
   assign A_chi[0][1][55]     = A[1][0][55] ^ ((~A[2][0][55]) & A[3][0][55]);
   assign A_chi[0][1][56]     = A[1][0][56] ^ ((~A[2][0][56]) & A[3][0][56]);
   assign A_chi[0][1][57]     = A[1][0][57] ^ ((~A[2][0][57]) & A[3][0][57]);
   assign A_chi[0][1][58]     = A[1][0][58] ^ ((~A[2][0][58]) & A[3][0][58]);
   assign A_chi[0][1][59]     = A[1][0][59] ^ ((~A[2][0][59]) & A[3][0][59]);
   assign A_chi[0][1][60]     = A[1][0][60] ^ ((~A[2][0][60]) & A[3][0][60]);
   assign A_chi[0][1][61]     = A[1][0][61] ^ ((~A[2][0][61]) & A[3][0][61]);
   assign A_chi[0][1][62]     = A[1][0][62] ^ ((~A[2][0][62]) & A[3][0][62]);
   assign A_chi[0][1][63]     = A[1][0][63] ^ ((~A[2][0][63]) & A[3][0][63]);
   assign A_chi[0][2][0]     = A[2][0][0] ^ ((~A[3][0][0]) & A[4][0][0]);
   assign A_chi[0][2][1]     = A[2][0][1] ^ ((~A[3][0][1]) & A[4][0][1]);
   assign A_chi[0][2][2]     = A[2][0][2] ^ ((~A[3][0][2]) & A[4][0][2]);
   assign A_chi[0][2][3]     = A[2][0][3] ^ ((~A[3][0][3]) & A[4][0][3]);
   assign A_chi[0][2][4]     = A[2][0][4] ^ ((~A[3][0][4]) & A[4][0][4]);
   assign A_chi[0][2][5]     = A[2][0][5] ^ ((~A[3][0][5]) & A[4][0][5]);
   assign A_chi[0][2][6]     = A[2][0][6] ^ ((~A[3][0][6]) & A[4][0][6]);
   assign A_chi[0][2][7]     = A[2][0][7] ^ ((~A[3][0][7]) & A[4][0][7]);
   assign A_chi[0][2][8]     = A[2][0][8] ^ ((~A[3][0][8]) & A[4][0][8]);
   assign A_chi[0][2][9]     = A[2][0][9] ^ ((~A[3][0][9]) & A[4][0][9]);
   assign A_chi[0][2][10]     = A[2][0][10] ^ ((~A[3][0][10]) & A[4][0][10]);
   assign A_chi[0][2][11]     = A[2][0][11] ^ ((~A[3][0][11]) & A[4][0][11]);
   assign A_chi[0][2][12]     = A[2][0][12] ^ ((~A[3][0][12]) & A[4][0][12]);
   assign A_chi[0][2][13]     = A[2][0][13] ^ ((~A[3][0][13]) & A[4][0][13]);
   assign A_chi[0][2][14]     = A[2][0][14] ^ ((~A[3][0][14]) & A[4][0][14]);
   assign A_chi[0][2][15]     = A[2][0][15] ^ ((~A[3][0][15]) & A[4][0][15]);
   assign A_chi[0][2][16]     = A[2][0][16] ^ ((~A[3][0][16]) & A[4][0][16]);
   assign A_chi[0][2][17]     = A[2][0][17] ^ ((~A[3][0][17]) & A[4][0][17]);
   assign A_chi[0][2][18]     = A[2][0][18] ^ ((~A[3][0][18]) & A[4][0][18]);
   assign A_chi[0][2][19]     = A[2][0][19] ^ ((~A[3][0][19]) & A[4][0][19]);
   assign A_chi[0][2][20]     = A[2][0][20] ^ ((~A[3][0][20]) & A[4][0][20]);
   assign A_chi[0][2][21]     = A[2][0][21] ^ ((~A[3][0][21]) & A[4][0][21]);
   assign A_chi[0][2][22]     = A[2][0][22] ^ ((~A[3][0][22]) & A[4][0][22]);
   assign A_chi[0][2][23]     = A[2][0][23] ^ ((~A[3][0][23]) & A[4][0][23]);
   assign A_chi[0][2][24]     = A[2][0][24] ^ ((~A[3][0][24]) & A[4][0][24]);
   assign A_chi[0][2][25]     = A[2][0][25] ^ ((~A[3][0][25]) & A[4][0][25]);
   assign A_chi[0][2][26]     = A[2][0][26] ^ ((~A[3][0][26]) & A[4][0][26]);
   assign A_chi[0][2][27]     = A[2][0][27] ^ ((~A[3][0][27]) & A[4][0][27]);
   assign A_chi[0][2][28]     = A[2][0][28] ^ ((~A[3][0][28]) & A[4][0][28]);
   assign A_chi[0][2][29]     = A[2][0][29] ^ ((~A[3][0][29]) & A[4][0][29]);
   assign A_chi[0][2][30]     = A[2][0][30] ^ ((~A[3][0][30]) & A[4][0][30]);
   assign A_chi[0][2][31]     = A[2][0][31] ^ ((~A[3][0][31]) & A[4][0][31]);
   assign A_chi[0][2][32]     = A[2][0][32] ^ ((~A[3][0][32]) & A[4][0][32]);
   assign A_chi[0][2][33]     = A[2][0][33] ^ ((~A[3][0][33]) & A[4][0][33]);
   assign A_chi[0][2][34]     = A[2][0][34] ^ ((~A[3][0][34]) & A[4][0][34]);
   assign A_chi[0][2][35]     = A[2][0][35] ^ ((~A[3][0][35]) & A[4][0][35]);
   assign A_chi[0][2][36]     = A[2][0][36] ^ ((~A[3][0][36]) & A[4][0][36]);
   assign A_chi[0][2][37]     = A[2][0][37] ^ ((~A[3][0][37]) & A[4][0][37]);
   assign A_chi[0][2][38]     = A[2][0][38] ^ ((~A[3][0][38]) & A[4][0][38]);
   assign A_chi[0][2][39]     = A[2][0][39] ^ ((~A[3][0][39]) & A[4][0][39]);
   assign A_chi[0][2][40]     = A[2][0][40] ^ ((~A[3][0][40]) & A[4][0][40]);
   assign A_chi[0][2][41]     = A[2][0][41] ^ ((~A[3][0][41]) & A[4][0][41]);
   assign A_chi[0][2][42]     = A[2][0][42] ^ ((~A[3][0][42]) & A[4][0][42]);
   assign A_chi[0][2][43]     = A[2][0][43] ^ ((~A[3][0][43]) & A[4][0][43]);
   assign A_chi[0][2][44]     = A[2][0][44] ^ ((~A[3][0][44]) & A[4][0][44]);
   assign A_chi[0][2][45]     = A[2][0][45] ^ ((~A[3][0][45]) & A[4][0][45]);
   assign A_chi[0][2][46]     = A[2][0][46] ^ ((~A[3][0][46]) & A[4][0][46]);
   assign A_chi[0][2][47]     = A[2][0][47] ^ ((~A[3][0][47]) & A[4][0][47]);
   assign A_chi[0][2][48]     = A[2][0][48] ^ ((~A[3][0][48]) & A[4][0][48]);
   assign A_chi[0][2][49]     = A[2][0][49] ^ ((~A[3][0][49]) & A[4][0][49]);
   assign A_chi[0][2][50]     = A[2][0][50] ^ ((~A[3][0][50]) & A[4][0][50]);
   assign A_chi[0][2][51]     = A[2][0][51] ^ ((~A[3][0][51]) & A[4][0][51]);
   assign A_chi[0][2][52]     = A[2][0][52] ^ ((~A[3][0][52]) & A[4][0][52]);
   assign A_chi[0][2][53]     = A[2][0][53] ^ ((~A[3][0][53]) & A[4][0][53]);
   assign A_chi[0][2][54]     = A[2][0][54] ^ ((~A[3][0][54]) & A[4][0][54]);
   assign A_chi[0][2][55]     = A[2][0][55] ^ ((~A[3][0][55]) & A[4][0][55]);
   assign A_chi[0][2][56]     = A[2][0][56] ^ ((~A[3][0][56]) & A[4][0][56]);
   assign A_chi[0][2][57]     = A[2][0][57] ^ ((~A[3][0][57]) & A[4][0][57]);
   assign A_chi[0][2][58]     = A[2][0][58] ^ ((~A[3][0][58]) & A[4][0][58]);
   assign A_chi[0][2][59]     = A[2][0][59] ^ ((~A[3][0][59]) & A[4][0][59]);
   assign A_chi[0][2][60]     = A[2][0][60] ^ ((~A[3][0][60]) & A[4][0][60]);
   assign A_chi[0][2][61]     = A[2][0][61] ^ ((~A[3][0][61]) & A[4][0][61]);
   assign A_chi[0][2][62]     = A[2][0][62] ^ ((~A[3][0][62]) & A[4][0][62]);
   assign A_chi[0][2][63]     = A[2][0][63] ^ ((~A[3][0][63]) & A[4][0][63]);
   assign A_chi[0][3][0]     = A[3][0][0] ^ ((~A[4][0][0]) & A[0][0][0]);
   assign A_chi[0][3][1]     = A[3][0][1] ^ ((~A[4][0][1]) & A[0][0][1]);
   assign A_chi[0][3][2]     = A[3][0][2] ^ ((~A[4][0][2]) & A[0][0][2]);
   assign A_chi[0][3][3]     = A[3][0][3] ^ ((~A[4][0][3]) & A[0][0][3]);
   assign A_chi[0][3][4]     = A[3][0][4] ^ ((~A[4][0][4]) & A[0][0][4]);
   assign A_chi[0][3][5]     = A[3][0][5] ^ ((~A[4][0][5]) & A[0][0][5]);
   assign A_chi[0][3][6]     = A[3][0][6] ^ ((~A[4][0][6]) & A[0][0][6]);
   assign A_chi[0][3][7]     = A[3][0][7] ^ ((~A[4][0][7]) & A[0][0][7]);
   assign A_chi[0][3][8]     = A[3][0][8] ^ ((~A[4][0][8]) & A[0][0][8]);
   assign A_chi[0][3][9]     = A[3][0][9] ^ ((~A[4][0][9]) & A[0][0][9]);
   assign A_chi[0][3][10]     = A[3][0][10] ^ ((~A[4][0][10]) & A[0][0][10]);
   assign A_chi[0][3][11]     = A[3][0][11] ^ ((~A[4][0][11]) & A[0][0][11]);
   assign A_chi[0][3][12]     = A[3][0][12] ^ ((~A[4][0][12]) & A[0][0][12]);
   assign A_chi[0][3][13]     = A[3][0][13] ^ ((~A[4][0][13]) & A[0][0][13]);
   assign A_chi[0][3][14]     = A[3][0][14] ^ ((~A[4][0][14]) & A[0][0][14]);
   assign A_chi[0][3][15]     = A[3][0][15] ^ ((~A[4][0][15]) & A[0][0][15]);
   assign A_chi[0][3][16]     = A[3][0][16] ^ ((~A[4][0][16]) & A[0][0][16]);
   assign A_chi[0][3][17]     = A[3][0][17] ^ ((~A[4][0][17]) & A[0][0][17]);
   assign A_chi[0][3][18]     = A[3][0][18] ^ ((~A[4][0][18]) & A[0][0][18]);
   assign A_chi[0][3][19]     = A[3][0][19] ^ ((~A[4][0][19]) & A[0][0][19]);
   assign A_chi[0][3][20]     = A[3][0][20] ^ ((~A[4][0][20]) & A[0][0][20]);
   assign A_chi[0][3][21]     = A[3][0][21] ^ ((~A[4][0][21]) & A[0][0][21]);
   assign A_chi[0][3][22]     = A[3][0][22] ^ ((~A[4][0][22]) & A[0][0][22]);
   assign A_chi[0][3][23]     = A[3][0][23] ^ ((~A[4][0][23]) & A[0][0][23]);
   assign A_chi[0][3][24]     = A[3][0][24] ^ ((~A[4][0][24]) & A[0][0][24]);
   assign A_chi[0][3][25]     = A[3][0][25] ^ ((~A[4][0][25]) & A[0][0][25]);
   assign A_chi[0][3][26]     = A[3][0][26] ^ ((~A[4][0][26]) & A[0][0][26]);
   assign A_chi[0][3][27]     = A[3][0][27] ^ ((~A[4][0][27]) & A[0][0][27]);
   assign A_chi[0][3][28]     = A[3][0][28] ^ ((~A[4][0][28]) & A[0][0][28]);
   assign A_chi[0][3][29]     = A[3][0][29] ^ ((~A[4][0][29]) & A[0][0][29]);
   assign A_chi[0][3][30]     = A[3][0][30] ^ ((~A[4][0][30]) & A[0][0][30]);
   assign A_chi[0][3][31]     = A[3][0][31] ^ ((~A[4][0][31]) & A[0][0][31]);
   assign A_chi[0][3][32]     = A[3][0][32] ^ ((~A[4][0][32]) & A[0][0][32]);
   assign A_chi[0][3][33]     = A[3][0][33] ^ ((~A[4][0][33]) & A[0][0][33]);
   assign A_chi[0][3][34]     = A[3][0][34] ^ ((~A[4][0][34]) & A[0][0][34]);
   assign A_chi[0][3][35]     = A[3][0][35] ^ ((~A[4][0][35]) & A[0][0][35]);
   assign A_chi[0][3][36]     = A[3][0][36] ^ ((~A[4][0][36]) & A[0][0][36]);
   assign A_chi[0][3][37]     = A[3][0][37] ^ ((~A[4][0][37]) & A[0][0][37]);
   assign A_chi[0][3][38]     = A[3][0][38] ^ ((~A[4][0][38]) & A[0][0][38]);
   assign A_chi[0][3][39]     = A[3][0][39] ^ ((~A[4][0][39]) & A[0][0][39]);
   assign A_chi[0][3][40]     = A[3][0][40] ^ ((~A[4][0][40]) & A[0][0][40]);
   assign A_chi[0][3][41]     = A[3][0][41] ^ ((~A[4][0][41]) & A[0][0][41]);
   assign A_chi[0][3][42]     = A[3][0][42] ^ ((~A[4][0][42]) & A[0][0][42]);
   assign A_chi[0][3][43]     = A[3][0][43] ^ ((~A[4][0][43]) & A[0][0][43]);
   assign A_chi[0][3][44]     = A[3][0][44] ^ ((~A[4][0][44]) & A[0][0][44]);
   assign A_chi[0][3][45]     = A[3][0][45] ^ ((~A[4][0][45]) & A[0][0][45]);
   assign A_chi[0][3][46]     = A[3][0][46] ^ ((~A[4][0][46]) & A[0][0][46]);
   assign A_chi[0][3][47]     = A[3][0][47] ^ ((~A[4][0][47]) & A[0][0][47]);
   assign A_chi[0][3][48]     = A[3][0][48] ^ ((~A[4][0][48]) & A[0][0][48]);
   assign A_chi[0][3][49]     = A[3][0][49] ^ ((~A[4][0][49]) & A[0][0][49]);
   assign A_chi[0][3][50]     = A[3][0][50] ^ ((~A[4][0][50]) & A[0][0][50]);
   assign A_chi[0][3][51]     = A[3][0][51] ^ ((~A[4][0][51]) & A[0][0][51]);
   assign A_chi[0][3][52]     = A[3][0][52] ^ ((~A[4][0][52]) & A[0][0][52]);
   assign A_chi[0][3][53]     = A[3][0][53] ^ ((~A[4][0][53]) & A[0][0][53]);
   assign A_chi[0][3][54]     = A[3][0][54] ^ ((~A[4][0][54]) & A[0][0][54]);
   assign A_chi[0][3][55]     = A[3][0][55] ^ ((~A[4][0][55]) & A[0][0][55]);
   assign A_chi[0][3][56]     = A[3][0][56] ^ ((~A[4][0][56]) & A[0][0][56]);
   assign A_chi[0][3][57]     = A[3][0][57] ^ ((~A[4][0][57]) & A[0][0][57]);
   assign A_chi[0][3][58]     = A[3][0][58] ^ ((~A[4][0][58]) & A[0][0][58]);
   assign A_chi[0][3][59]     = A[3][0][59] ^ ((~A[4][0][59]) & A[0][0][59]);
   assign A_chi[0][3][60]     = A[3][0][60] ^ ((~A[4][0][60]) & A[0][0][60]);
   assign A_chi[0][3][61]     = A[3][0][61] ^ ((~A[4][0][61]) & A[0][0][61]);
   assign A_chi[0][3][62]     = A[3][0][62] ^ ((~A[4][0][62]) & A[0][0][62]);
   assign A_chi[0][3][63]     = A[3][0][63] ^ ((~A[4][0][63]) & A[0][0][63]);
   assign A_chi[0][4][0]     = A[4][0][0] ^ ((~A[0][0][0]) & A[1][0][0]);
   assign A_chi[0][4][1]     = A[4][0][1] ^ ((~A[0][0][1]) & A[1][0][1]);
   assign A_chi[0][4][2]     = A[4][0][2] ^ ((~A[0][0][2]) & A[1][0][2]);
   assign A_chi[0][4][3]     = A[4][0][3] ^ ((~A[0][0][3]) & A[1][0][3]);
   assign A_chi[0][4][4]     = A[4][0][4] ^ ((~A[0][0][4]) & A[1][0][4]);
   assign A_chi[0][4][5]     = A[4][0][5] ^ ((~A[0][0][5]) & A[1][0][5]);
   assign A_chi[0][4][6]     = A[4][0][6] ^ ((~A[0][0][6]) & A[1][0][6]);
   assign A_chi[0][4][7]     = A[4][0][7] ^ ((~A[0][0][7]) & A[1][0][7]);
   assign A_chi[0][4][8]     = A[4][0][8] ^ ((~A[0][0][8]) & A[1][0][8]);
   assign A_chi[0][4][9]     = A[4][0][9] ^ ((~A[0][0][9]) & A[1][0][9]);
   assign A_chi[0][4][10]     = A[4][0][10] ^ ((~A[0][0][10]) & A[1][0][10]);
   assign A_chi[0][4][11]     = A[4][0][11] ^ ((~A[0][0][11]) & A[1][0][11]);
   assign A_chi[0][4][12]     = A[4][0][12] ^ ((~A[0][0][12]) & A[1][0][12]);
   assign A_chi[0][4][13]     = A[4][0][13] ^ ((~A[0][0][13]) & A[1][0][13]);
   assign A_chi[0][4][14]     = A[4][0][14] ^ ((~A[0][0][14]) & A[1][0][14]);
   assign A_chi[0][4][15]     = A[4][0][15] ^ ((~A[0][0][15]) & A[1][0][15]);
   assign A_chi[0][4][16]     = A[4][0][16] ^ ((~A[0][0][16]) & A[1][0][16]);
   assign A_chi[0][4][17]     = A[4][0][17] ^ ((~A[0][0][17]) & A[1][0][17]);
   assign A_chi[0][4][18]     = A[4][0][18] ^ ((~A[0][0][18]) & A[1][0][18]);
   assign A_chi[0][4][19]     = A[4][0][19] ^ ((~A[0][0][19]) & A[1][0][19]);
   assign A_chi[0][4][20]     = A[4][0][20] ^ ((~A[0][0][20]) & A[1][0][20]);
   assign A_chi[0][4][21]     = A[4][0][21] ^ ((~A[0][0][21]) & A[1][0][21]);
   assign A_chi[0][4][22]     = A[4][0][22] ^ ((~A[0][0][22]) & A[1][0][22]);
   assign A_chi[0][4][23]     = A[4][0][23] ^ ((~A[0][0][23]) & A[1][0][23]);
   assign A_chi[0][4][24]     = A[4][0][24] ^ ((~A[0][0][24]) & A[1][0][24]);
   assign A_chi[0][4][25]     = A[4][0][25] ^ ((~A[0][0][25]) & A[1][0][25]);
   assign A_chi[0][4][26]     = A[4][0][26] ^ ((~A[0][0][26]) & A[1][0][26]);
   assign A_chi[0][4][27]     = A[4][0][27] ^ ((~A[0][0][27]) & A[1][0][27]);
   assign A_chi[0][4][28]     = A[4][0][28] ^ ((~A[0][0][28]) & A[1][0][28]);
   assign A_chi[0][4][29]     = A[4][0][29] ^ ((~A[0][0][29]) & A[1][0][29]);
   assign A_chi[0][4][30]     = A[4][0][30] ^ ((~A[0][0][30]) & A[1][0][30]);
   assign A_chi[0][4][31]     = A[4][0][31] ^ ((~A[0][0][31]) & A[1][0][31]);
   assign A_chi[0][4][32]     = A[4][0][32] ^ ((~A[0][0][32]) & A[1][0][32]);
   assign A_chi[0][4][33]     = A[4][0][33] ^ ((~A[0][0][33]) & A[1][0][33]);
   assign A_chi[0][4][34]     = A[4][0][34] ^ ((~A[0][0][34]) & A[1][0][34]);
   assign A_chi[0][4][35]     = A[4][0][35] ^ ((~A[0][0][35]) & A[1][0][35]);
   assign A_chi[0][4][36]     = A[4][0][36] ^ ((~A[0][0][36]) & A[1][0][36]);
   assign A_chi[0][4][37]     = A[4][0][37] ^ ((~A[0][0][37]) & A[1][0][37]);
   assign A_chi[0][4][38]     = A[4][0][38] ^ ((~A[0][0][38]) & A[1][0][38]);
   assign A_chi[0][4][39]     = A[4][0][39] ^ ((~A[0][0][39]) & A[1][0][39]);
   assign A_chi[0][4][40]     = A[4][0][40] ^ ((~A[0][0][40]) & A[1][0][40]);
   assign A_chi[0][4][41]     = A[4][0][41] ^ ((~A[0][0][41]) & A[1][0][41]);
   assign A_chi[0][4][42]     = A[4][0][42] ^ ((~A[0][0][42]) & A[1][0][42]);
   assign A_chi[0][4][43]     = A[4][0][43] ^ ((~A[0][0][43]) & A[1][0][43]);
   assign A_chi[0][4][44]     = A[4][0][44] ^ ((~A[0][0][44]) & A[1][0][44]);
   assign A_chi[0][4][45]     = A[4][0][45] ^ ((~A[0][0][45]) & A[1][0][45]);
   assign A_chi[0][4][46]     = A[4][0][46] ^ ((~A[0][0][46]) & A[1][0][46]);
   assign A_chi[0][4][47]     = A[4][0][47] ^ ((~A[0][0][47]) & A[1][0][47]);
   assign A_chi[0][4][48]     = A[4][0][48] ^ ((~A[0][0][48]) & A[1][0][48]);
   assign A_chi[0][4][49]     = A[4][0][49] ^ ((~A[0][0][49]) & A[1][0][49]);
   assign A_chi[0][4][50]     = A[4][0][50] ^ ((~A[0][0][50]) & A[1][0][50]);
   assign A_chi[0][4][51]     = A[4][0][51] ^ ((~A[0][0][51]) & A[1][0][51]);
   assign A_chi[0][4][52]     = A[4][0][52] ^ ((~A[0][0][52]) & A[1][0][52]);
   assign A_chi[0][4][53]     = A[4][0][53] ^ ((~A[0][0][53]) & A[1][0][53]);
   assign A_chi[0][4][54]     = A[4][0][54] ^ ((~A[0][0][54]) & A[1][0][54]);
   assign A_chi[0][4][55]     = A[4][0][55] ^ ((~A[0][0][55]) & A[1][0][55]);
   assign A_chi[0][4][56]     = A[4][0][56] ^ ((~A[0][0][56]) & A[1][0][56]);
   assign A_chi[0][4][57]     = A[4][0][57] ^ ((~A[0][0][57]) & A[1][0][57]);
   assign A_chi[0][4][58]     = A[4][0][58] ^ ((~A[0][0][58]) & A[1][0][58]);
   assign A_chi[0][4][59]     = A[4][0][59] ^ ((~A[0][0][59]) & A[1][0][59]);
   assign A_chi[0][4][60]     = A[4][0][60] ^ ((~A[0][0][60]) & A[1][0][60]);
   assign A_chi[0][4][61]     = A[4][0][61] ^ ((~A[0][0][61]) & A[1][0][61]);
   assign A_chi[0][4][62]     = A[4][0][62] ^ ((~A[0][0][62]) & A[1][0][62]);
   assign A_chi[0][4][63]     = A[4][0][63] ^ ((~A[0][0][63]) & A[1][0][63]);
   assign A_chi[1][0][0]     = A[0][1][0] ^ ((~A[1][1][0]) & A[2][1][0]);
   assign A_chi[1][0][1]     = A[0][1][1] ^ ((~A[1][1][1]) & A[2][1][1]);
   assign A_chi[1][0][2]     = A[0][1][2] ^ ((~A[1][1][2]) & A[2][1][2]);
   assign A_chi[1][0][3]     = A[0][1][3] ^ ((~A[1][1][3]) & A[2][1][3]);
   assign A_chi[1][0][4]     = A[0][1][4] ^ ((~A[1][1][4]) & A[2][1][4]);
   assign A_chi[1][0][5]     = A[0][1][5] ^ ((~A[1][1][5]) & A[2][1][5]);
   assign A_chi[1][0][6]     = A[0][1][6] ^ ((~A[1][1][6]) & A[2][1][6]);
   assign A_chi[1][0][7]     = A[0][1][7] ^ ((~A[1][1][7]) & A[2][1][7]);
   assign A_chi[1][0][8]     = A[0][1][8] ^ ((~A[1][1][8]) & A[2][1][8]);
   assign A_chi[1][0][9]     = A[0][1][9] ^ ((~A[1][1][9]) & A[2][1][9]);
   assign A_chi[1][0][10]     = A[0][1][10] ^ ((~A[1][1][10]) & A[2][1][10]);
   assign A_chi[1][0][11]     = A[0][1][11] ^ ((~A[1][1][11]) & A[2][1][11]);
   assign A_chi[1][0][12]     = A[0][1][12] ^ ((~A[1][1][12]) & A[2][1][12]);
   assign A_chi[1][0][13]     = A[0][1][13] ^ ((~A[1][1][13]) & A[2][1][13]);
   assign A_chi[1][0][14]     = A[0][1][14] ^ ((~A[1][1][14]) & A[2][1][14]);
   assign A_chi[1][0][15]     = A[0][1][15] ^ ((~A[1][1][15]) & A[2][1][15]);
   assign A_chi[1][0][16]     = A[0][1][16] ^ ((~A[1][1][16]) & A[2][1][16]);
   assign A_chi[1][0][17]     = A[0][1][17] ^ ((~A[1][1][17]) & A[2][1][17]);
   assign A_chi[1][0][18]     = A[0][1][18] ^ ((~A[1][1][18]) & A[2][1][18]);
   assign A_chi[1][0][19]     = A[0][1][19] ^ ((~A[1][1][19]) & A[2][1][19]);
   assign A_chi[1][0][20]     = A[0][1][20] ^ ((~A[1][1][20]) & A[2][1][20]);
   assign A_chi[1][0][21]     = A[0][1][21] ^ ((~A[1][1][21]) & A[2][1][21]);
   assign A_chi[1][0][22]     = A[0][1][22] ^ ((~A[1][1][22]) & A[2][1][22]);
   assign A_chi[1][0][23]     = A[0][1][23] ^ ((~A[1][1][23]) & A[2][1][23]);
   assign A_chi[1][0][24]     = A[0][1][24] ^ ((~A[1][1][24]) & A[2][1][24]);
   assign A_chi[1][0][25]     = A[0][1][25] ^ ((~A[1][1][25]) & A[2][1][25]);
   assign A_chi[1][0][26]     = A[0][1][26] ^ ((~A[1][1][26]) & A[2][1][26]);
   assign A_chi[1][0][27]     = A[0][1][27] ^ ((~A[1][1][27]) & A[2][1][27]);
   assign A_chi[1][0][28]     = A[0][1][28] ^ ((~A[1][1][28]) & A[2][1][28]);
   assign A_chi[1][0][29]     = A[0][1][29] ^ ((~A[1][1][29]) & A[2][1][29]);
   assign A_chi[1][0][30]     = A[0][1][30] ^ ((~A[1][1][30]) & A[2][1][30]);
   assign A_chi[1][0][31]     = A[0][1][31] ^ ((~A[1][1][31]) & A[2][1][31]);
   assign A_chi[1][0][32]     = A[0][1][32] ^ ((~A[1][1][32]) & A[2][1][32]);
   assign A_chi[1][0][33]     = A[0][1][33] ^ ((~A[1][1][33]) & A[2][1][33]);
   assign A_chi[1][0][34]     = A[0][1][34] ^ ((~A[1][1][34]) & A[2][1][34]);
   assign A_chi[1][0][35]     = A[0][1][35] ^ ((~A[1][1][35]) & A[2][1][35]);
   assign A_chi[1][0][36]     = A[0][1][36] ^ ((~A[1][1][36]) & A[2][1][36]);
   assign A_chi[1][0][37]     = A[0][1][37] ^ ((~A[1][1][37]) & A[2][1][37]);
   assign A_chi[1][0][38]     = A[0][1][38] ^ ((~A[1][1][38]) & A[2][1][38]);
   assign A_chi[1][0][39]     = A[0][1][39] ^ ((~A[1][1][39]) & A[2][1][39]);
   assign A_chi[1][0][40]     = A[0][1][40] ^ ((~A[1][1][40]) & A[2][1][40]);
   assign A_chi[1][0][41]     = A[0][1][41] ^ ((~A[1][1][41]) & A[2][1][41]);
   assign A_chi[1][0][42]     = A[0][1][42] ^ ((~A[1][1][42]) & A[2][1][42]);
   assign A_chi[1][0][43]     = A[0][1][43] ^ ((~A[1][1][43]) & A[2][1][43]);
   assign A_chi[1][0][44]     = A[0][1][44] ^ ((~A[1][1][44]) & A[2][1][44]);
   assign A_chi[1][0][45]     = A[0][1][45] ^ ((~A[1][1][45]) & A[2][1][45]);
   assign A_chi[1][0][46]     = A[0][1][46] ^ ((~A[1][1][46]) & A[2][1][46]);
   assign A_chi[1][0][47]     = A[0][1][47] ^ ((~A[1][1][47]) & A[2][1][47]);
   assign A_chi[1][0][48]     = A[0][1][48] ^ ((~A[1][1][48]) & A[2][1][48]);
   assign A_chi[1][0][49]     = A[0][1][49] ^ ((~A[1][1][49]) & A[2][1][49]);
   assign A_chi[1][0][50]     = A[0][1][50] ^ ((~A[1][1][50]) & A[2][1][50]);
   assign A_chi[1][0][51]     = A[0][1][51] ^ ((~A[1][1][51]) & A[2][1][51]);
   assign A_chi[1][0][52]     = A[0][1][52] ^ ((~A[1][1][52]) & A[2][1][52]);
   assign A_chi[1][0][53]     = A[0][1][53] ^ ((~A[1][1][53]) & A[2][1][53]);
   assign A_chi[1][0][54]     = A[0][1][54] ^ ((~A[1][1][54]) & A[2][1][54]);
   assign A_chi[1][0][55]     = A[0][1][55] ^ ((~A[1][1][55]) & A[2][1][55]);
   assign A_chi[1][0][56]     = A[0][1][56] ^ ((~A[1][1][56]) & A[2][1][56]);
   assign A_chi[1][0][57]     = A[0][1][57] ^ ((~A[1][1][57]) & A[2][1][57]);
   assign A_chi[1][0][58]     = A[0][1][58] ^ ((~A[1][1][58]) & A[2][1][58]);
   assign A_chi[1][0][59]     = A[0][1][59] ^ ((~A[1][1][59]) & A[2][1][59]);
   assign A_chi[1][0][60]     = A[0][1][60] ^ ((~A[1][1][60]) & A[2][1][60]);
   assign A_chi[1][0][61]     = A[0][1][61] ^ ((~A[1][1][61]) & A[2][1][61]);
   assign A_chi[1][0][62]     = A[0][1][62] ^ ((~A[1][1][62]) & A[2][1][62]);
   assign A_chi[1][0][63]     = A[0][1][63] ^ ((~A[1][1][63]) & A[2][1][63]);
   assign A_chi[1][1][0]     = A[1][1][0] ^ ((~A[2][1][0]) & A[3][1][0]);
   assign A_chi[1][1][1]     = A[1][1][1] ^ ((~A[2][1][1]) & A[3][1][1]);
   assign A_chi[1][1][2]     = A[1][1][2] ^ ((~A[2][1][2]) & A[3][1][2]);
   assign A_chi[1][1][3]     = A[1][1][3] ^ ((~A[2][1][3]) & A[3][1][3]);
   assign A_chi[1][1][4]     = A[1][1][4] ^ ((~A[2][1][4]) & A[3][1][4]);
   assign A_chi[1][1][5]     = A[1][1][5] ^ ((~A[2][1][5]) & A[3][1][5]);
   assign A_chi[1][1][6]     = A[1][1][6] ^ ((~A[2][1][6]) & A[3][1][6]);
   assign A_chi[1][1][7]     = A[1][1][7] ^ ((~A[2][1][7]) & A[3][1][7]);
   assign A_chi[1][1][8]     = A[1][1][8] ^ ((~A[2][1][8]) & A[3][1][8]);
   assign A_chi[1][1][9]     = A[1][1][9] ^ ((~A[2][1][9]) & A[3][1][9]);
   assign A_chi[1][1][10]     = A[1][1][10] ^ ((~A[2][1][10]) & A[3][1][10]);
   assign A_chi[1][1][11]     = A[1][1][11] ^ ((~A[2][1][11]) & A[3][1][11]);
   assign A_chi[1][1][12]     = A[1][1][12] ^ ((~A[2][1][12]) & A[3][1][12]);
   assign A_chi[1][1][13]     = A[1][1][13] ^ ((~A[2][1][13]) & A[3][1][13]);
   assign A_chi[1][1][14]     = A[1][1][14] ^ ((~A[2][1][14]) & A[3][1][14]);
   assign A_chi[1][1][15]     = A[1][1][15] ^ ((~A[2][1][15]) & A[3][1][15]);
   assign A_chi[1][1][16]     = A[1][1][16] ^ ((~A[2][1][16]) & A[3][1][16]);
   assign A_chi[1][1][17]     = A[1][1][17] ^ ((~A[2][1][17]) & A[3][1][17]);
   assign A_chi[1][1][18]     = A[1][1][18] ^ ((~A[2][1][18]) & A[3][1][18]);
   assign A_chi[1][1][19]     = A[1][1][19] ^ ((~A[2][1][19]) & A[3][1][19]);
   assign A_chi[1][1][20]     = A[1][1][20] ^ ((~A[2][1][20]) & A[3][1][20]);
   assign A_chi[1][1][21]     = A[1][1][21] ^ ((~A[2][1][21]) & A[3][1][21]);
   assign A_chi[1][1][22]     = A[1][1][22] ^ ((~A[2][1][22]) & A[3][1][22]);
   assign A_chi[1][1][23]     = A[1][1][23] ^ ((~A[2][1][23]) & A[3][1][23]);
   assign A_chi[1][1][24]     = A[1][1][24] ^ ((~A[2][1][24]) & A[3][1][24]);
   assign A_chi[1][1][25]     = A[1][1][25] ^ ((~A[2][1][25]) & A[3][1][25]);
   assign A_chi[1][1][26]     = A[1][1][26] ^ ((~A[2][1][26]) & A[3][1][26]);
   assign A_chi[1][1][27]     = A[1][1][27] ^ ((~A[2][1][27]) & A[3][1][27]);
   assign A_chi[1][1][28]     = A[1][1][28] ^ ((~A[2][1][28]) & A[3][1][28]);
   assign A_chi[1][1][29]     = A[1][1][29] ^ ((~A[2][1][29]) & A[3][1][29]);
   assign A_chi[1][1][30]     = A[1][1][30] ^ ((~A[2][1][30]) & A[3][1][30]);
   assign A_chi[1][1][31]     = A[1][1][31] ^ ((~A[2][1][31]) & A[3][1][31]);
   assign A_chi[1][1][32]     = A[1][1][32] ^ ((~A[2][1][32]) & A[3][1][32]);
   assign A_chi[1][1][33]     = A[1][1][33] ^ ((~A[2][1][33]) & A[3][1][33]);
   assign A_chi[1][1][34]     = A[1][1][34] ^ ((~A[2][1][34]) & A[3][1][34]);
   assign A_chi[1][1][35]     = A[1][1][35] ^ ((~A[2][1][35]) & A[3][1][35]);
   assign A_chi[1][1][36]     = A[1][1][36] ^ ((~A[2][1][36]) & A[3][1][36]);
   assign A_chi[1][1][37]     = A[1][1][37] ^ ((~A[2][1][37]) & A[3][1][37]);
   assign A_chi[1][1][38]     = A[1][1][38] ^ ((~A[2][1][38]) & A[3][1][38]);
   assign A_chi[1][1][39]     = A[1][1][39] ^ ((~A[2][1][39]) & A[3][1][39]);
   assign A_chi[1][1][40]     = A[1][1][40] ^ ((~A[2][1][40]) & A[3][1][40]);
   assign A_chi[1][1][41]     = A[1][1][41] ^ ((~A[2][1][41]) & A[3][1][41]);
   assign A_chi[1][1][42]     = A[1][1][42] ^ ((~A[2][1][42]) & A[3][1][42]);
   assign A_chi[1][1][43]     = A[1][1][43] ^ ((~A[2][1][43]) & A[3][1][43]);
   assign A_chi[1][1][44]     = A[1][1][44] ^ ((~A[2][1][44]) & A[3][1][44]);
   assign A_chi[1][1][45]     = A[1][1][45] ^ ((~A[2][1][45]) & A[3][1][45]);
   assign A_chi[1][1][46]     = A[1][1][46] ^ ((~A[2][1][46]) & A[3][1][46]);
   assign A_chi[1][1][47]     = A[1][1][47] ^ ((~A[2][1][47]) & A[3][1][47]);
   assign A_chi[1][1][48]     = A[1][1][48] ^ ((~A[2][1][48]) & A[3][1][48]);
   assign A_chi[1][1][49]     = A[1][1][49] ^ ((~A[2][1][49]) & A[3][1][49]);
   assign A_chi[1][1][50]     = A[1][1][50] ^ ((~A[2][1][50]) & A[3][1][50]);
   assign A_chi[1][1][51]     = A[1][1][51] ^ ((~A[2][1][51]) & A[3][1][51]);
   assign A_chi[1][1][52]     = A[1][1][52] ^ ((~A[2][1][52]) & A[3][1][52]);
   assign A_chi[1][1][53]     = A[1][1][53] ^ ((~A[2][1][53]) & A[3][1][53]);
   assign A_chi[1][1][54]     = A[1][1][54] ^ ((~A[2][1][54]) & A[3][1][54]);
   assign A_chi[1][1][55]     = A[1][1][55] ^ ((~A[2][1][55]) & A[3][1][55]);
   assign A_chi[1][1][56]     = A[1][1][56] ^ ((~A[2][1][56]) & A[3][1][56]);
   assign A_chi[1][1][57]     = A[1][1][57] ^ ((~A[2][1][57]) & A[3][1][57]);
   assign A_chi[1][1][58]     = A[1][1][58] ^ ((~A[2][1][58]) & A[3][1][58]);
   assign A_chi[1][1][59]     = A[1][1][59] ^ ((~A[2][1][59]) & A[3][1][59]);
   assign A_chi[1][1][60]     = A[1][1][60] ^ ((~A[2][1][60]) & A[3][1][60]);
   assign A_chi[1][1][61]     = A[1][1][61] ^ ((~A[2][1][61]) & A[3][1][61]);
   assign A_chi[1][1][62]     = A[1][1][62] ^ ((~A[2][1][62]) & A[3][1][62]);
   assign A_chi[1][1][63]     = A[1][1][63] ^ ((~A[2][1][63]) & A[3][1][63]);
   assign A_chi[1][2][0]     = A[2][1][0] ^ ((~A[3][1][0]) & A[4][1][0]);
   assign A_chi[1][2][1]     = A[2][1][1] ^ ((~A[3][1][1]) & A[4][1][1]);
   assign A_chi[1][2][2]     = A[2][1][2] ^ ((~A[3][1][2]) & A[4][1][2]);
   assign A_chi[1][2][3]     = A[2][1][3] ^ ((~A[3][1][3]) & A[4][1][3]);
   assign A_chi[1][2][4]     = A[2][1][4] ^ ((~A[3][1][4]) & A[4][1][4]);
   assign A_chi[1][2][5]     = A[2][1][5] ^ ((~A[3][1][5]) & A[4][1][5]);
   assign A_chi[1][2][6]     = A[2][1][6] ^ ((~A[3][1][6]) & A[4][1][6]);
   assign A_chi[1][2][7]     = A[2][1][7] ^ ((~A[3][1][7]) & A[4][1][7]);
   assign A_chi[1][2][8]     = A[2][1][8] ^ ((~A[3][1][8]) & A[4][1][8]);
   assign A_chi[1][2][9]     = A[2][1][9] ^ ((~A[3][1][9]) & A[4][1][9]);
   assign A_chi[1][2][10]     = A[2][1][10] ^ ((~A[3][1][10]) & A[4][1][10]);
   assign A_chi[1][2][11]     = A[2][1][11] ^ ((~A[3][1][11]) & A[4][1][11]);
   assign A_chi[1][2][12]     = A[2][1][12] ^ ((~A[3][1][12]) & A[4][1][12]);
   assign A_chi[1][2][13]     = A[2][1][13] ^ ((~A[3][1][13]) & A[4][1][13]);
   assign A_chi[1][2][14]     = A[2][1][14] ^ ((~A[3][1][14]) & A[4][1][14]);
   assign A_chi[1][2][15]     = A[2][1][15] ^ ((~A[3][1][15]) & A[4][1][15]);
   assign A_chi[1][2][16]     = A[2][1][16] ^ ((~A[3][1][16]) & A[4][1][16]);
   assign A_chi[1][2][17]     = A[2][1][17] ^ ((~A[3][1][17]) & A[4][1][17]);
   assign A_chi[1][2][18]     = A[2][1][18] ^ ((~A[3][1][18]) & A[4][1][18]);
   assign A_chi[1][2][19]     = A[2][1][19] ^ ((~A[3][1][19]) & A[4][1][19]);
   assign A_chi[1][2][20]     = A[2][1][20] ^ ((~A[3][1][20]) & A[4][1][20]);
   assign A_chi[1][2][21]     = A[2][1][21] ^ ((~A[3][1][21]) & A[4][1][21]);
   assign A_chi[1][2][22]     = A[2][1][22] ^ ((~A[3][1][22]) & A[4][1][22]);
   assign A_chi[1][2][23]     = A[2][1][23] ^ ((~A[3][1][23]) & A[4][1][23]);
   assign A_chi[1][2][24]     = A[2][1][24] ^ ((~A[3][1][24]) & A[4][1][24]);
   assign A_chi[1][2][25]     = A[2][1][25] ^ ((~A[3][1][25]) & A[4][1][25]);
   assign A_chi[1][2][26]     = A[2][1][26] ^ ((~A[3][1][26]) & A[4][1][26]);
   assign A_chi[1][2][27]     = A[2][1][27] ^ ((~A[3][1][27]) & A[4][1][27]);
   assign A_chi[1][2][28]     = A[2][1][28] ^ ((~A[3][1][28]) & A[4][1][28]);
   assign A_chi[1][2][29]     = A[2][1][29] ^ ((~A[3][1][29]) & A[4][1][29]);
   assign A_chi[1][2][30]     = A[2][1][30] ^ ((~A[3][1][30]) & A[4][1][30]);
   assign A_chi[1][2][31]     = A[2][1][31] ^ ((~A[3][1][31]) & A[4][1][31]);
   assign A_chi[1][2][32]     = A[2][1][32] ^ ((~A[3][1][32]) & A[4][1][32]);
   assign A_chi[1][2][33]     = A[2][1][33] ^ ((~A[3][1][33]) & A[4][1][33]);
   assign A_chi[1][2][34]     = A[2][1][34] ^ ((~A[3][1][34]) & A[4][1][34]);
   assign A_chi[1][2][35]     = A[2][1][35] ^ ((~A[3][1][35]) & A[4][1][35]);
   assign A_chi[1][2][36]     = A[2][1][36] ^ ((~A[3][1][36]) & A[4][1][36]);
   assign A_chi[1][2][37]     = A[2][1][37] ^ ((~A[3][1][37]) & A[4][1][37]);
   assign A_chi[1][2][38]     = A[2][1][38] ^ ((~A[3][1][38]) & A[4][1][38]);
   assign A_chi[1][2][39]     = A[2][1][39] ^ ((~A[3][1][39]) & A[4][1][39]);
   assign A_chi[1][2][40]     = A[2][1][40] ^ ((~A[3][1][40]) & A[4][1][40]);
   assign A_chi[1][2][41]     = A[2][1][41] ^ ((~A[3][1][41]) & A[4][1][41]);
   assign A_chi[1][2][42]     = A[2][1][42] ^ ((~A[3][1][42]) & A[4][1][42]);
   assign A_chi[1][2][43]     = A[2][1][43] ^ ((~A[3][1][43]) & A[4][1][43]);
   assign A_chi[1][2][44]     = A[2][1][44] ^ ((~A[3][1][44]) & A[4][1][44]);
   assign A_chi[1][2][45]     = A[2][1][45] ^ ((~A[3][1][45]) & A[4][1][45]);
   assign A_chi[1][2][46]     = A[2][1][46] ^ ((~A[3][1][46]) & A[4][1][46]);
   assign A_chi[1][2][47]     = A[2][1][47] ^ ((~A[3][1][47]) & A[4][1][47]);
   assign A_chi[1][2][48]     = A[2][1][48] ^ ((~A[3][1][48]) & A[4][1][48]);
   assign A_chi[1][2][49]     = A[2][1][49] ^ ((~A[3][1][49]) & A[4][1][49]);
   assign A_chi[1][2][50]     = A[2][1][50] ^ ((~A[3][1][50]) & A[4][1][50]);
   assign A_chi[1][2][51]     = A[2][1][51] ^ ((~A[3][1][51]) & A[4][1][51]);
   assign A_chi[1][2][52]     = A[2][1][52] ^ ((~A[3][1][52]) & A[4][1][52]);
   assign A_chi[1][2][53]     = A[2][1][53] ^ ((~A[3][1][53]) & A[4][1][53]);
   assign A_chi[1][2][54]     = A[2][1][54] ^ ((~A[3][1][54]) & A[4][1][54]);
   assign A_chi[1][2][55]     = A[2][1][55] ^ ((~A[3][1][55]) & A[4][1][55]);
   assign A_chi[1][2][56]     = A[2][1][56] ^ ((~A[3][1][56]) & A[4][1][56]);
   assign A_chi[1][2][57]     = A[2][1][57] ^ ((~A[3][1][57]) & A[4][1][57]);
   assign A_chi[1][2][58]     = A[2][1][58] ^ ((~A[3][1][58]) & A[4][1][58]);
   assign A_chi[1][2][59]     = A[2][1][59] ^ ((~A[3][1][59]) & A[4][1][59]);
   assign A_chi[1][2][60]     = A[2][1][60] ^ ((~A[3][1][60]) & A[4][1][60]);
   assign A_chi[1][2][61]     = A[2][1][61] ^ ((~A[3][1][61]) & A[4][1][61]);
   assign A_chi[1][2][62]     = A[2][1][62] ^ ((~A[3][1][62]) & A[4][1][62]);
   assign A_chi[1][2][63]     = A[2][1][63] ^ ((~A[3][1][63]) & A[4][1][63]);
   assign A_chi[1][3][0]     = A[3][1][0] ^ ((~A[4][1][0]) & A[0][1][0]);
   assign A_chi[1][3][1]     = A[3][1][1] ^ ((~A[4][1][1]) & A[0][1][1]);
   assign A_chi[1][3][2]     = A[3][1][2] ^ ((~A[4][1][2]) & A[0][1][2]);
   assign A_chi[1][3][3]     = A[3][1][3] ^ ((~A[4][1][3]) & A[0][1][3]);
   assign A_chi[1][3][4]     = A[3][1][4] ^ ((~A[4][1][4]) & A[0][1][4]);
   assign A_chi[1][3][5]     = A[3][1][5] ^ ((~A[4][1][5]) & A[0][1][5]);
   assign A_chi[1][3][6]     = A[3][1][6] ^ ((~A[4][1][6]) & A[0][1][6]);
   assign A_chi[1][3][7]     = A[3][1][7] ^ ((~A[4][1][7]) & A[0][1][7]);
   assign A_chi[1][3][8]     = A[3][1][8] ^ ((~A[4][1][8]) & A[0][1][8]);
   assign A_chi[1][3][9]     = A[3][1][9] ^ ((~A[4][1][9]) & A[0][1][9]);
   assign A_chi[1][3][10]     = A[3][1][10] ^ ((~A[4][1][10]) & A[0][1][10]);
   assign A_chi[1][3][11]     = A[3][1][11] ^ ((~A[4][1][11]) & A[0][1][11]);
   assign A_chi[1][3][12]     = A[3][1][12] ^ ((~A[4][1][12]) & A[0][1][12]);
   assign A_chi[1][3][13]     = A[3][1][13] ^ ((~A[4][1][13]) & A[0][1][13]);
   assign A_chi[1][3][14]     = A[3][1][14] ^ ((~A[4][1][14]) & A[0][1][14]);
   assign A_chi[1][3][15]     = A[3][1][15] ^ ((~A[4][1][15]) & A[0][1][15]);
   assign A_chi[1][3][16]     = A[3][1][16] ^ ((~A[4][1][16]) & A[0][1][16]);
   assign A_chi[1][3][17]     = A[3][1][17] ^ ((~A[4][1][17]) & A[0][1][17]);
   assign A_chi[1][3][18]     = A[3][1][18] ^ ((~A[4][1][18]) & A[0][1][18]);
   assign A_chi[1][3][19]     = A[3][1][19] ^ ((~A[4][1][19]) & A[0][1][19]);
   assign A_chi[1][3][20]     = A[3][1][20] ^ ((~A[4][1][20]) & A[0][1][20]);
   assign A_chi[1][3][21]     = A[3][1][21] ^ ((~A[4][1][21]) & A[0][1][21]);
   assign A_chi[1][3][22]     = A[3][1][22] ^ ((~A[4][1][22]) & A[0][1][22]);
   assign A_chi[1][3][23]     = A[3][1][23] ^ ((~A[4][1][23]) & A[0][1][23]);
   assign A_chi[1][3][24]     = A[3][1][24] ^ ((~A[4][1][24]) & A[0][1][24]);
   assign A_chi[1][3][25]     = A[3][1][25] ^ ((~A[4][1][25]) & A[0][1][25]);
   assign A_chi[1][3][26]     = A[3][1][26] ^ ((~A[4][1][26]) & A[0][1][26]);
   assign A_chi[1][3][27]     = A[3][1][27] ^ ((~A[4][1][27]) & A[0][1][27]);
   assign A_chi[1][3][28]     = A[3][1][28] ^ ((~A[4][1][28]) & A[0][1][28]);
   assign A_chi[1][3][29]     = A[3][1][29] ^ ((~A[4][1][29]) & A[0][1][29]);
   assign A_chi[1][3][30]     = A[3][1][30] ^ ((~A[4][1][30]) & A[0][1][30]);
   assign A_chi[1][3][31]     = A[3][1][31] ^ ((~A[4][1][31]) & A[0][1][31]);
   assign A_chi[1][3][32]     = A[3][1][32] ^ ((~A[4][1][32]) & A[0][1][32]);
   assign A_chi[1][3][33]     = A[3][1][33] ^ ((~A[4][1][33]) & A[0][1][33]);
   assign A_chi[1][3][34]     = A[3][1][34] ^ ((~A[4][1][34]) & A[0][1][34]);
   assign A_chi[1][3][35]     = A[3][1][35] ^ ((~A[4][1][35]) & A[0][1][35]);
   assign A_chi[1][3][36]     = A[3][1][36] ^ ((~A[4][1][36]) & A[0][1][36]);
   assign A_chi[1][3][37]     = A[3][1][37] ^ ((~A[4][1][37]) & A[0][1][37]);
   assign A_chi[1][3][38]     = A[3][1][38] ^ ((~A[4][1][38]) & A[0][1][38]);
   assign A_chi[1][3][39]     = A[3][1][39] ^ ((~A[4][1][39]) & A[0][1][39]);
   assign A_chi[1][3][40]     = A[3][1][40] ^ ((~A[4][1][40]) & A[0][1][40]);
   assign A_chi[1][3][41]     = A[3][1][41] ^ ((~A[4][1][41]) & A[0][1][41]);
   assign A_chi[1][3][42]     = A[3][1][42] ^ ((~A[4][1][42]) & A[0][1][42]);
   assign A_chi[1][3][43]     = A[3][1][43] ^ ((~A[4][1][43]) & A[0][1][43]);
   assign A_chi[1][3][44]     = A[3][1][44] ^ ((~A[4][1][44]) & A[0][1][44]);
   assign A_chi[1][3][45]     = A[3][1][45] ^ ((~A[4][1][45]) & A[0][1][45]);
   assign A_chi[1][3][46]     = A[3][1][46] ^ ((~A[4][1][46]) & A[0][1][46]);
   assign A_chi[1][3][47]     = A[3][1][47] ^ ((~A[4][1][47]) & A[0][1][47]);
   assign A_chi[1][3][48]     = A[3][1][48] ^ ((~A[4][1][48]) & A[0][1][48]);
   assign A_chi[1][3][49]     = A[3][1][49] ^ ((~A[4][1][49]) & A[0][1][49]);
   assign A_chi[1][3][50]     = A[3][1][50] ^ ((~A[4][1][50]) & A[0][1][50]);
   assign A_chi[1][3][51]     = A[3][1][51] ^ ((~A[4][1][51]) & A[0][1][51]);
   assign A_chi[1][3][52]     = A[3][1][52] ^ ((~A[4][1][52]) & A[0][1][52]);
   assign A_chi[1][3][53]     = A[3][1][53] ^ ((~A[4][1][53]) & A[0][1][53]);
   assign A_chi[1][3][54]     = A[3][1][54] ^ ((~A[4][1][54]) & A[0][1][54]);
   assign A_chi[1][3][55]     = A[3][1][55] ^ ((~A[4][1][55]) & A[0][1][55]);
   assign A_chi[1][3][56]     = A[3][1][56] ^ ((~A[4][1][56]) & A[0][1][56]);
   assign A_chi[1][3][57]     = A[3][1][57] ^ ((~A[4][1][57]) & A[0][1][57]);
   assign A_chi[1][3][58]     = A[3][1][58] ^ ((~A[4][1][58]) & A[0][1][58]);
   assign A_chi[1][3][59]     = A[3][1][59] ^ ((~A[4][1][59]) & A[0][1][59]);
   assign A_chi[1][3][60]     = A[3][1][60] ^ ((~A[4][1][60]) & A[0][1][60]);
   assign A_chi[1][3][61]     = A[3][1][61] ^ ((~A[4][1][61]) & A[0][1][61]);
   assign A_chi[1][3][62]     = A[3][1][62] ^ ((~A[4][1][62]) & A[0][1][62]);
   assign A_chi[1][3][63]     = A[3][1][63] ^ ((~A[4][1][63]) & A[0][1][63]);
   assign A_chi[1][4][0]     = A[4][1][0] ^ ((~A[0][1][0]) & A[1][1][0]);
   assign A_chi[1][4][1]     = A[4][1][1] ^ ((~A[0][1][1]) & A[1][1][1]);
   assign A_chi[1][4][2]     = A[4][1][2] ^ ((~A[0][1][2]) & A[1][1][2]);
   assign A_chi[1][4][3]     = A[4][1][3] ^ ((~A[0][1][3]) & A[1][1][3]);
   assign A_chi[1][4][4]     = A[4][1][4] ^ ((~A[0][1][4]) & A[1][1][4]);
   assign A_chi[1][4][5]     = A[4][1][5] ^ ((~A[0][1][5]) & A[1][1][5]);
   assign A_chi[1][4][6]     = A[4][1][6] ^ ((~A[0][1][6]) & A[1][1][6]);
   assign A_chi[1][4][7]     = A[4][1][7] ^ ((~A[0][1][7]) & A[1][1][7]);
   assign A_chi[1][4][8]     = A[4][1][8] ^ ((~A[0][1][8]) & A[1][1][8]);
   assign A_chi[1][4][9]     = A[4][1][9] ^ ((~A[0][1][9]) & A[1][1][9]);
   assign A_chi[1][4][10]     = A[4][1][10] ^ ((~A[0][1][10]) & A[1][1][10]);
   assign A_chi[1][4][11]     = A[4][1][11] ^ ((~A[0][1][11]) & A[1][1][11]);
   assign A_chi[1][4][12]     = A[4][1][12] ^ ((~A[0][1][12]) & A[1][1][12]);
   assign A_chi[1][4][13]     = A[4][1][13] ^ ((~A[0][1][13]) & A[1][1][13]);
   assign A_chi[1][4][14]     = A[4][1][14] ^ ((~A[0][1][14]) & A[1][1][14]);
   assign A_chi[1][4][15]     = A[4][1][15] ^ ((~A[0][1][15]) & A[1][1][15]);
   assign A_chi[1][4][16]     = A[4][1][16] ^ ((~A[0][1][16]) & A[1][1][16]);
   assign A_chi[1][4][17]     = A[4][1][17] ^ ((~A[0][1][17]) & A[1][1][17]);
   assign A_chi[1][4][18]     = A[4][1][18] ^ ((~A[0][1][18]) & A[1][1][18]);
   assign A_chi[1][4][19]     = A[4][1][19] ^ ((~A[0][1][19]) & A[1][1][19]);
   assign A_chi[1][4][20]     = A[4][1][20] ^ ((~A[0][1][20]) & A[1][1][20]);
   assign A_chi[1][4][21]     = A[4][1][21] ^ ((~A[0][1][21]) & A[1][1][21]);
   assign A_chi[1][4][22]     = A[4][1][22] ^ ((~A[0][1][22]) & A[1][1][22]);
   assign A_chi[1][4][23]     = A[4][1][23] ^ ((~A[0][1][23]) & A[1][1][23]);
   assign A_chi[1][4][24]     = A[4][1][24] ^ ((~A[0][1][24]) & A[1][1][24]);
   assign A_chi[1][4][25]     = A[4][1][25] ^ ((~A[0][1][25]) & A[1][1][25]);
   assign A_chi[1][4][26]     = A[4][1][26] ^ ((~A[0][1][26]) & A[1][1][26]);
   assign A_chi[1][4][27]     = A[4][1][27] ^ ((~A[0][1][27]) & A[1][1][27]);
   assign A_chi[1][4][28]     = A[4][1][28] ^ ((~A[0][1][28]) & A[1][1][28]);
   assign A_chi[1][4][29]     = A[4][1][29] ^ ((~A[0][1][29]) & A[1][1][29]);
   assign A_chi[1][4][30]     = A[4][1][30] ^ ((~A[0][1][30]) & A[1][1][30]);
   assign A_chi[1][4][31]     = A[4][1][31] ^ ((~A[0][1][31]) & A[1][1][31]);
   assign A_chi[1][4][32]     = A[4][1][32] ^ ((~A[0][1][32]) & A[1][1][32]);
   assign A_chi[1][4][33]     = A[4][1][33] ^ ((~A[0][1][33]) & A[1][1][33]);
   assign A_chi[1][4][34]     = A[4][1][34] ^ ((~A[0][1][34]) & A[1][1][34]);
   assign A_chi[1][4][35]     = A[4][1][35] ^ ((~A[0][1][35]) & A[1][1][35]);
   assign A_chi[1][4][36]     = A[4][1][36] ^ ((~A[0][1][36]) & A[1][1][36]);
   assign A_chi[1][4][37]     = A[4][1][37] ^ ((~A[0][1][37]) & A[1][1][37]);
   assign A_chi[1][4][38]     = A[4][1][38] ^ ((~A[0][1][38]) & A[1][1][38]);
   assign A_chi[1][4][39]     = A[4][1][39] ^ ((~A[0][1][39]) & A[1][1][39]);
   assign A_chi[1][4][40]     = A[4][1][40] ^ ((~A[0][1][40]) & A[1][1][40]);
   assign A_chi[1][4][41]     = A[4][1][41] ^ ((~A[0][1][41]) & A[1][1][41]);
   assign A_chi[1][4][42]     = A[4][1][42] ^ ((~A[0][1][42]) & A[1][1][42]);
   assign A_chi[1][4][43]     = A[4][1][43] ^ ((~A[0][1][43]) & A[1][1][43]);
   assign A_chi[1][4][44]     = A[4][1][44] ^ ((~A[0][1][44]) & A[1][1][44]);
   assign A_chi[1][4][45]     = A[4][1][45] ^ ((~A[0][1][45]) & A[1][1][45]);
   assign A_chi[1][4][46]     = A[4][1][46] ^ ((~A[0][1][46]) & A[1][1][46]);
   assign A_chi[1][4][47]     = A[4][1][47] ^ ((~A[0][1][47]) & A[1][1][47]);
   assign A_chi[1][4][48]     = A[4][1][48] ^ ((~A[0][1][48]) & A[1][1][48]);
   assign A_chi[1][4][49]     = A[4][1][49] ^ ((~A[0][1][49]) & A[1][1][49]);
   assign A_chi[1][4][50]     = A[4][1][50] ^ ((~A[0][1][50]) & A[1][1][50]);
   assign A_chi[1][4][51]     = A[4][1][51] ^ ((~A[0][1][51]) & A[1][1][51]);
   assign A_chi[1][4][52]     = A[4][1][52] ^ ((~A[0][1][52]) & A[1][1][52]);
   assign A_chi[1][4][53]     = A[4][1][53] ^ ((~A[0][1][53]) & A[1][1][53]);
   assign A_chi[1][4][54]     = A[4][1][54] ^ ((~A[0][1][54]) & A[1][1][54]);
   assign A_chi[1][4][55]     = A[4][1][55] ^ ((~A[0][1][55]) & A[1][1][55]);
   assign A_chi[1][4][56]     = A[4][1][56] ^ ((~A[0][1][56]) & A[1][1][56]);
   assign A_chi[1][4][57]     = A[4][1][57] ^ ((~A[0][1][57]) & A[1][1][57]);
   assign A_chi[1][4][58]     = A[4][1][58] ^ ((~A[0][1][58]) & A[1][1][58]);
   assign A_chi[1][4][59]     = A[4][1][59] ^ ((~A[0][1][59]) & A[1][1][59]);
   assign A_chi[1][4][60]     = A[4][1][60] ^ ((~A[0][1][60]) & A[1][1][60]);
   assign A_chi[1][4][61]     = A[4][1][61] ^ ((~A[0][1][61]) & A[1][1][61]);
   assign A_chi[1][4][62]     = A[4][1][62] ^ ((~A[0][1][62]) & A[1][1][62]);
   assign A_chi[1][4][63]     = A[4][1][63] ^ ((~A[0][1][63]) & A[1][1][63]);
   assign A_chi[2][0][0]     = A[0][2][0] ^ ((~A[1][2][0]) & A[2][2][0]);
   assign A_chi[2][0][1]     = A[0][2][1] ^ ((~A[1][2][1]) & A[2][2][1]);
   assign A_chi[2][0][2]     = A[0][2][2] ^ ((~A[1][2][2]) & A[2][2][2]);
   assign A_chi[2][0][3]     = A[0][2][3] ^ ((~A[1][2][3]) & A[2][2][3]);
   assign A_chi[2][0][4]     = A[0][2][4] ^ ((~A[1][2][4]) & A[2][2][4]);
   assign A_chi[2][0][5]     = A[0][2][5] ^ ((~A[1][2][5]) & A[2][2][5]);
   assign A_chi[2][0][6]     = A[0][2][6] ^ ((~A[1][2][6]) & A[2][2][6]);
   assign A_chi[2][0][7]     = A[0][2][7] ^ ((~A[1][2][7]) & A[2][2][7]);
   assign A_chi[2][0][8]     = A[0][2][8] ^ ((~A[1][2][8]) & A[2][2][8]);
   assign A_chi[2][0][9]     = A[0][2][9] ^ ((~A[1][2][9]) & A[2][2][9]);
   assign A_chi[2][0][10]     = A[0][2][10] ^ ((~A[1][2][10]) & A[2][2][10]);
   assign A_chi[2][0][11]     = A[0][2][11] ^ ((~A[1][2][11]) & A[2][2][11]);
   assign A_chi[2][0][12]     = A[0][2][12] ^ ((~A[1][2][12]) & A[2][2][12]);
   assign A_chi[2][0][13]     = A[0][2][13] ^ ((~A[1][2][13]) & A[2][2][13]);
   assign A_chi[2][0][14]     = A[0][2][14] ^ ((~A[1][2][14]) & A[2][2][14]);
   assign A_chi[2][0][15]     = A[0][2][15] ^ ((~A[1][2][15]) & A[2][2][15]);
   assign A_chi[2][0][16]     = A[0][2][16] ^ ((~A[1][2][16]) & A[2][2][16]);
   assign A_chi[2][0][17]     = A[0][2][17] ^ ((~A[1][2][17]) & A[2][2][17]);
   assign A_chi[2][0][18]     = A[0][2][18] ^ ((~A[1][2][18]) & A[2][2][18]);
   assign A_chi[2][0][19]     = A[0][2][19] ^ ((~A[1][2][19]) & A[2][2][19]);
   assign A_chi[2][0][20]     = A[0][2][20] ^ ((~A[1][2][20]) & A[2][2][20]);
   assign A_chi[2][0][21]     = A[0][2][21] ^ ((~A[1][2][21]) & A[2][2][21]);
   assign A_chi[2][0][22]     = A[0][2][22] ^ ((~A[1][2][22]) & A[2][2][22]);
   assign A_chi[2][0][23]     = A[0][2][23] ^ ((~A[1][2][23]) & A[2][2][23]);
   assign A_chi[2][0][24]     = A[0][2][24] ^ ((~A[1][2][24]) & A[2][2][24]);
   assign A_chi[2][0][25]     = A[0][2][25] ^ ((~A[1][2][25]) & A[2][2][25]);
   assign A_chi[2][0][26]     = A[0][2][26] ^ ((~A[1][2][26]) & A[2][2][26]);
   assign A_chi[2][0][27]     = A[0][2][27] ^ ((~A[1][2][27]) & A[2][2][27]);
   assign A_chi[2][0][28]     = A[0][2][28] ^ ((~A[1][2][28]) & A[2][2][28]);
   assign A_chi[2][0][29]     = A[0][2][29] ^ ((~A[1][2][29]) & A[2][2][29]);
   assign A_chi[2][0][30]     = A[0][2][30] ^ ((~A[1][2][30]) & A[2][2][30]);
   assign A_chi[2][0][31]     = A[0][2][31] ^ ((~A[1][2][31]) & A[2][2][31]);
   assign A_chi[2][0][32]     = A[0][2][32] ^ ((~A[1][2][32]) & A[2][2][32]);
   assign A_chi[2][0][33]     = A[0][2][33] ^ ((~A[1][2][33]) & A[2][2][33]);
   assign A_chi[2][0][34]     = A[0][2][34] ^ ((~A[1][2][34]) & A[2][2][34]);
   assign A_chi[2][0][35]     = A[0][2][35] ^ ((~A[1][2][35]) & A[2][2][35]);
   assign A_chi[2][0][36]     = A[0][2][36] ^ ((~A[1][2][36]) & A[2][2][36]);
   assign A_chi[2][0][37]     = A[0][2][37] ^ ((~A[1][2][37]) & A[2][2][37]);
   assign A_chi[2][0][38]     = A[0][2][38] ^ ((~A[1][2][38]) & A[2][2][38]);
   assign A_chi[2][0][39]     = A[0][2][39] ^ ((~A[1][2][39]) & A[2][2][39]);
   assign A_chi[2][0][40]     = A[0][2][40] ^ ((~A[1][2][40]) & A[2][2][40]);
   assign A_chi[2][0][41]     = A[0][2][41] ^ ((~A[1][2][41]) & A[2][2][41]);
   assign A_chi[2][0][42]     = A[0][2][42] ^ ((~A[1][2][42]) & A[2][2][42]);
   assign A_chi[2][0][43]     = A[0][2][43] ^ ((~A[1][2][43]) & A[2][2][43]);
   assign A_chi[2][0][44]     = A[0][2][44] ^ ((~A[1][2][44]) & A[2][2][44]);
   assign A_chi[2][0][45]     = A[0][2][45] ^ ((~A[1][2][45]) & A[2][2][45]);
   assign A_chi[2][0][46]     = A[0][2][46] ^ ((~A[1][2][46]) & A[2][2][46]);
   assign A_chi[2][0][47]     = A[0][2][47] ^ ((~A[1][2][47]) & A[2][2][47]);
   assign A_chi[2][0][48]     = A[0][2][48] ^ ((~A[1][2][48]) & A[2][2][48]);
   assign A_chi[2][0][49]     = A[0][2][49] ^ ((~A[1][2][49]) & A[2][2][49]);
   assign A_chi[2][0][50]     = A[0][2][50] ^ ((~A[1][2][50]) & A[2][2][50]);
   assign A_chi[2][0][51]     = A[0][2][51] ^ ((~A[1][2][51]) & A[2][2][51]);
   assign A_chi[2][0][52]     = A[0][2][52] ^ ((~A[1][2][52]) & A[2][2][52]);
   assign A_chi[2][0][53]     = A[0][2][53] ^ ((~A[1][2][53]) & A[2][2][53]);
   assign A_chi[2][0][54]     = A[0][2][54] ^ ((~A[1][2][54]) & A[2][2][54]);
   assign A_chi[2][0][55]     = A[0][2][55] ^ ((~A[1][2][55]) & A[2][2][55]);
   assign A_chi[2][0][56]     = A[0][2][56] ^ ((~A[1][2][56]) & A[2][2][56]);
   assign A_chi[2][0][57]     = A[0][2][57] ^ ((~A[1][2][57]) & A[2][2][57]);
   assign A_chi[2][0][58]     = A[0][2][58] ^ ((~A[1][2][58]) & A[2][2][58]);
   assign A_chi[2][0][59]     = A[0][2][59] ^ ((~A[1][2][59]) & A[2][2][59]);
   assign A_chi[2][0][60]     = A[0][2][60] ^ ((~A[1][2][60]) & A[2][2][60]);
   assign A_chi[2][0][61]     = A[0][2][61] ^ ((~A[1][2][61]) & A[2][2][61]);
   assign A_chi[2][0][62]     = A[0][2][62] ^ ((~A[1][2][62]) & A[2][2][62]);
   assign A_chi[2][0][63]     = A[0][2][63] ^ ((~A[1][2][63]) & A[2][2][63]);
   assign A_chi[2][1][0]     = A[1][2][0] ^ ((~A[2][2][0]) & A[3][2][0]);
   assign A_chi[2][1][1]     = A[1][2][1] ^ ((~A[2][2][1]) & A[3][2][1]);
   assign A_chi[2][1][2]     = A[1][2][2] ^ ((~A[2][2][2]) & A[3][2][2]);
   assign A_chi[2][1][3]     = A[1][2][3] ^ ((~A[2][2][3]) & A[3][2][3]);
   assign A_chi[2][1][4]     = A[1][2][4] ^ ((~A[2][2][4]) & A[3][2][4]);
   assign A_chi[2][1][5]     = A[1][2][5] ^ ((~A[2][2][5]) & A[3][2][5]);
   assign A_chi[2][1][6]     = A[1][2][6] ^ ((~A[2][2][6]) & A[3][2][6]);
   assign A_chi[2][1][7]     = A[1][2][7] ^ ((~A[2][2][7]) & A[3][2][7]);
   assign A_chi[2][1][8]     = A[1][2][8] ^ ((~A[2][2][8]) & A[3][2][8]);
   assign A_chi[2][1][9]     = A[1][2][9] ^ ((~A[2][2][9]) & A[3][2][9]);
   assign A_chi[2][1][10]     = A[1][2][10] ^ ((~A[2][2][10]) & A[3][2][10]);
   assign A_chi[2][1][11]     = A[1][2][11] ^ ((~A[2][2][11]) & A[3][2][11]);
   assign A_chi[2][1][12]     = A[1][2][12] ^ ((~A[2][2][12]) & A[3][2][12]);
   assign A_chi[2][1][13]     = A[1][2][13] ^ ((~A[2][2][13]) & A[3][2][13]);
   assign A_chi[2][1][14]     = A[1][2][14] ^ ((~A[2][2][14]) & A[3][2][14]);
   assign A_chi[2][1][15]     = A[1][2][15] ^ ((~A[2][2][15]) & A[3][2][15]);
   assign A_chi[2][1][16]     = A[1][2][16] ^ ((~A[2][2][16]) & A[3][2][16]);
   assign A_chi[2][1][17]     = A[1][2][17] ^ ((~A[2][2][17]) & A[3][2][17]);
   assign A_chi[2][1][18]     = A[1][2][18] ^ ((~A[2][2][18]) & A[3][2][18]);
   assign A_chi[2][1][19]     = A[1][2][19] ^ ((~A[2][2][19]) & A[3][2][19]);
   assign A_chi[2][1][20]     = A[1][2][20] ^ ((~A[2][2][20]) & A[3][2][20]);
   assign A_chi[2][1][21]     = A[1][2][21] ^ ((~A[2][2][21]) & A[3][2][21]);
   assign A_chi[2][1][22]     = A[1][2][22] ^ ((~A[2][2][22]) & A[3][2][22]);
   assign A_chi[2][1][23]     = A[1][2][23] ^ ((~A[2][2][23]) & A[3][2][23]);
   assign A_chi[2][1][24]     = A[1][2][24] ^ ((~A[2][2][24]) & A[3][2][24]);
   assign A_chi[2][1][25]     = A[1][2][25] ^ ((~A[2][2][25]) & A[3][2][25]);
   assign A_chi[2][1][26]     = A[1][2][26] ^ ((~A[2][2][26]) & A[3][2][26]);
   assign A_chi[2][1][27]     = A[1][2][27] ^ ((~A[2][2][27]) & A[3][2][27]);
   assign A_chi[2][1][28]     = A[1][2][28] ^ ((~A[2][2][28]) & A[3][2][28]);
   assign A_chi[2][1][29]     = A[1][2][29] ^ ((~A[2][2][29]) & A[3][2][29]);
   assign A_chi[2][1][30]     = A[1][2][30] ^ ((~A[2][2][30]) & A[3][2][30]);
   assign A_chi[2][1][31]     = A[1][2][31] ^ ((~A[2][2][31]) & A[3][2][31]);
   assign A_chi[2][1][32]     = A[1][2][32] ^ ((~A[2][2][32]) & A[3][2][32]);
   assign A_chi[2][1][33]     = A[1][2][33] ^ ((~A[2][2][33]) & A[3][2][33]);
   assign A_chi[2][1][34]     = A[1][2][34] ^ ((~A[2][2][34]) & A[3][2][34]);
   assign A_chi[2][1][35]     = A[1][2][35] ^ ((~A[2][2][35]) & A[3][2][35]);
   assign A_chi[2][1][36]     = A[1][2][36] ^ ((~A[2][2][36]) & A[3][2][36]);
   assign A_chi[2][1][37]     = A[1][2][37] ^ ((~A[2][2][37]) & A[3][2][37]);
   assign A_chi[2][1][38]     = A[1][2][38] ^ ((~A[2][2][38]) & A[3][2][38]);
   assign A_chi[2][1][39]     = A[1][2][39] ^ ((~A[2][2][39]) & A[3][2][39]);
   assign A_chi[2][1][40]     = A[1][2][40] ^ ((~A[2][2][40]) & A[3][2][40]);
   assign A_chi[2][1][41]     = A[1][2][41] ^ ((~A[2][2][41]) & A[3][2][41]);
   assign A_chi[2][1][42]     = A[1][2][42] ^ ((~A[2][2][42]) & A[3][2][42]);
   assign A_chi[2][1][43]     = A[1][2][43] ^ ((~A[2][2][43]) & A[3][2][43]);
   assign A_chi[2][1][44]     = A[1][2][44] ^ ((~A[2][2][44]) & A[3][2][44]);
   assign A_chi[2][1][45]     = A[1][2][45] ^ ((~A[2][2][45]) & A[3][2][45]);
   assign A_chi[2][1][46]     = A[1][2][46] ^ ((~A[2][2][46]) & A[3][2][46]);
   assign A_chi[2][1][47]     = A[1][2][47] ^ ((~A[2][2][47]) & A[3][2][47]);
   assign A_chi[2][1][48]     = A[1][2][48] ^ ((~A[2][2][48]) & A[3][2][48]);
   assign A_chi[2][1][49]     = A[1][2][49] ^ ((~A[2][2][49]) & A[3][2][49]);
   assign A_chi[2][1][50]     = A[1][2][50] ^ ((~A[2][2][50]) & A[3][2][50]);
   assign A_chi[2][1][51]     = A[1][2][51] ^ ((~A[2][2][51]) & A[3][2][51]);
   assign A_chi[2][1][52]     = A[1][2][52] ^ ((~A[2][2][52]) & A[3][2][52]);
   assign A_chi[2][1][53]     = A[1][2][53] ^ ((~A[2][2][53]) & A[3][2][53]);
   assign A_chi[2][1][54]     = A[1][2][54] ^ ((~A[2][2][54]) & A[3][2][54]);
   assign A_chi[2][1][55]     = A[1][2][55] ^ ((~A[2][2][55]) & A[3][2][55]);
   assign A_chi[2][1][56]     = A[1][2][56] ^ ((~A[2][2][56]) & A[3][2][56]);
   assign A_chi[2][1][57]     = A[1][2][57] ^ ((~A[2][2][57]) & A[3][2][57]);
   assign A_chi[2][1][58]     = A[1][2][58] ^ ((~A[2][2][58]) & A[3][2][58]);
   assign A_chi[2][1][59]     = A[1][2][59] ^ ((~A[2][2][59]) & A[3][2][59]);
   assign A_chi[2][1][60]     = A[1][2][60] ^ ((~A[2][2][60]) & A[3][2][60]);
   assign A_chi[2][1][61]     = A[1][2][61] ^ ((~A[2][2][61]) & A[3][2][61]);
   assign A_chi[2][1][62]     = A[1][2][62] ^ ((~A[2][2][62]) & A[3][2][62]);
   assign A_chi[2][1][63]     = A[1][2][63] ^ ((~A[2][2][63]) & A[3][2][63]);
   assign A_chi[2][2][0]     = A[2][2][0] ^ ((~A[3][2][0]) & A[4][2][0]);
   assign A_chi[2][2][1]     = A[2][2][1] ^ ((~A[3][2][1]) & A[4][2][1]);
   assign A_chi[2][2][2]     = A[2][2][2] ^ ((~A[3][2][2]) & A[4][2][2]);
   assign A_chi[2][2][3]     = A[2][2][3] ^ ((~A[3][2][3]) & A[4][2][3]);
   assign A_chi[2][2][4]     = A[2][2][4] ^ ((~A[3][2][4]) & A[4][2][4]);
   assign A_chi[2][2][5]     = A[2][2][5] ^ ((~A[3][2][5]) & A[4][2][5]);
   assign A_chi[2][2][6]     = A[2][2][6] ^ ((~A[3][2][6]) & A[4][2][6]);
   assign A_chi[2][2][7]     = A[2][2][7] ^ ((~A[3][2][7]) & A[4][2][7]);
   assign A_chi[2][2][8]     = A[2][2][8] ^ ((~A[3][2][8]) & A[4][2][8]);
   assign A_chi[2][2][9]     = A[2][2][9] ^ ((~A[3][2][9]) & A[4][2][9]);
   assign A_chi[2][2][10]     = A[2][2][10] ^ ((~A[3][2][10]) & A[4][2][10]);
   assign A_chi[2][2][11]     = A[2][2][11] ^ ((~A[3][2][11]) & A[4][2][11]);
   assign A_chi[2][2][12]     = A[2][2][12] ^ ((~A[3][2][12]) & A[4][2][12]);
   assign A_chi[2][2][13]     = A[2][2][13] ^ ((~A[3][2][13]) & A[4][2][13]);
   assign A_chi[2][2][14]     = A[2][2][14] ^ ((~A[3][2][14]) & A[4][2][14]);
   assign A_chi[2][2][15]     = A[2][2][15] ^ ((~A[3][2][15]) & A[4][2][15]);
   assign A_chi[2][2][16]     = A[2][2][16] ^ ((~A[3][2][16]) & A[4][2][16]);
   assign A_chi[2][2][17]     = A[2][2][17] ^ ((~A[3][2][17]) & A[4][2][17]);
   assign A_chi[2][2][18]     = A[2][2][18] ^ ((~A[3][2][18]) & A[4][2][18]);
   assign A_chi[2][2][19]     = A[2][2][19] ^ ((~A[3][2][19]) & A[4][2][19]);
   assign A_chi[2][2][20]     = A[2][2][20] ^ ((~A[3][2][20]) & A[4][2][20]);
   assign A_chi[2][2][21]     = A[2][2][21] ^ ((~A[3][2][21]) & A[4][2][21]);
   assign A_chi[2][2][22]     = A[2][2][22] ^ ((~A[3][2][22]) & A[4][2][22]);
   assign A_chi[2][2][23]     = A[2][2][23] ^ ((~A[3][2][23]) & A[4][2][23]);
   assign A_chi[2][2][24]     = A[2][2][24] ^ ((~A[3][2][24]) & A[4][2][24]);
   assign A_chi[2][2][25]     = A[2][2][25] ^ ((~A[3][2][25]) & A[4][2][25]);
   assign A_chi[2][2][26]     = A[2][2][26] ^ ((~A[3][2][26]) & A[4][2][26]);
   assign A_chi[2][2][27]     = A[2][2][27] ^ ((~A[3][2][27]) & A[4][2][27]);
   assign A_chi[2][2][28]     = A[2][2][28] ^ ((~A[3][2][28]) & A[4][2][28]);
   assign A_chi[2][2][29]     = A[2][2][29] ^ ((~A[3][2][29]) & A[4][2][29]);
   assign A_chi[2][2][30]     = A[2][2][30] ^ ((~A[3][2][30]) & A[4][2][30]);
   assign A_chi[2][2][31]     = A[2][2][31] ^ ((~A[3][2][31]) & A[4][2][31]);
   assign A_chi[2][2][32]     = A[2][2][32] ^ ((~A[3][2][32]) & A[4][2][32]);
   assign A_chi[2][2][33]     = A[2][2][33] ^ ((~A[3][2][33]) & A[4][2][33]);
   assign A_chi[2][2][34]     = A[2][2][34] ^ ((~A[3][2][34]) & A[4][2][34]);
   assign A_chi[2][2][35]     = A[2][2][35] ^ ((~A[3][2][35]) & A[4][2][35]);
   assign A_chi[2][2][36]     = A[2][2][36] ^ ((~A[3][2][36]) & A[4][2][36]);
   assign A_chi[2][2][37]     = A[2][2][37] ^ ((~A[3][2][37]) & A[4][2][37]);
   assign A_chi[2][2][38]     = A[2][2][38] ^ ((~A[3][2][38]) & A[4][2][38]);
   assign A_chi[2][2][39]     = A[2][2][39] ^ ((~A[3][2][39]) & A[4][2][39]);
   assign A_chi[2][2][40]     = A[2][2][40] ^ ((~A[3][2][40]) & A[4][2][40]);
   assign A_chi[2][2][41]     = A[2][2][41] ^ ((~A[3][2][41]) & A[4][2][41]);
   assign A_chi[2][2][42]     = A[2][2][42] ^ ((~A[3][2][42]) & A[4][2][42]);
   assign A_chi[2][2][43]     = A[2][2][43] ^ ((~A[3][2][43]) & A[4][2][43]);
   assign A_chi[2][2][44]     = A[2][2][44] ^ ((~A[3][2][44]) & A[4][2][44]);
   assign A_chi[2][2][45]     = A[2][2][45] ^ ((~A[3][2][45]) & A[4][2][45]);
   assign A_chi[2][2][46]     = A[2][2][46] ^ ((~A[3][2][46]) & A[4][2][46]);
   assign A_chi[2][2][47]     = A[2][2][47] ^ ((~A[3][2][47]) & A[4][2][47]);
   assign A_chi[2][2][48]     = A[2][2][48] ^ ((~A[3][2][48]) & A[4][2][48]);
   assign A_chi[2][2][49]     = A[2][2][49] ^ ((~A[3][2][49]) & A[4][2][49]);
   assign A_chi[2][2][50]     = A[2][2][50] ^ ((~A[3][2][50]) & A[4][2][50]);
   assign A_chi[2][2][51]     = A[2][2][51] ^ ((~A[3][2][51]) & A[4][2][51]);
   assign A_chi[2][2][52]     = A[2][2][52] ^ ((~A[3][2][52]) & A[4][2][52]);
   assign A_chi[2][2][53]     = A[2][2][53] ^ ((~A[3][2][53]) & A[4][2][53]);
   assign A_chi[2][2][54]     = A[2][2][54] ^ ((~A[3][2][54]) & A[4][2][54]);
   assign A_chi[2][2][55]     = A[2][2][55] ^ ((~A[3][2][55]) & A[4][2][55]);
   assign A_chi[2][2][56]     = A[2][2][56] ^ ((~A[3][2][56]) & A[4][2][56]);
   assign A_chi[2][2][57]     = A[2][2][57] ^ ((~A[3][2][57]) & A[4][2][57]);
   assign A_chi[2][2][58]     = A[2][2][58] ^ ((~A[3][2][58]) & A[4][2][58]);
   assign A_chi[2][2][59]     = A[2][2][59] ^ ((~A[3][2][59]) & A[4][2][59]);
   assign A_chi[2][2][60]     = A[2][2][60] ^ ((~A[3][2][60]) & A[4][2][60]);
   assign A_chi[2][2][61]     = A[2][2][61] ^ ((~A[3][2][61]) & A[4][2][61]);
   assign A_chi[2][2][62]     = A[2][2][62] ^ ((~A[3][2][62]) & A[4][2][62]);
   assign A_chi[2][2][63]     = A[2][2][63] ^ ((~A[3][2][63]) & A[4][2][63]);
   assign A_chi[2][3][0]     = A[3][2][0] ^ ((~A[4][2][0]) & A[0][2][0]);
   assign A_chi[2][3][1]     = A[3][2][1] ^ ((~A[4][2][1]) & A[0][2][1]);
   assign A_chi[2][3][2]     = A[3][2][2] ^ ((~A[4][2][2]) & A[0][2][2]);
   assign A_chi[2][3][3]     = A[3][2][3] ^ ((~A[4][2][3]) & A[0][2][3]);
   assign A_chi[2][3][4]     = A[3][2][4] ^ ((~A[4][2][4]) & A[0][2][4]);
   assign A_chi[2][3][5]     = A[3][2][5] ^ ((~A[4][2][5]) & A[0][2][5]);
   assign A_chi[2][3][6]     = A[3][2][6] ^ ((~A[4][2][6]) & A[0][2][6]);
   assign A_chi[2][3][7]     = A[3][2][7] ^ ((~A[4][2][7]) & A[0][2][7]);
   assign A_chi[2][3][8]     = A[3][2][8] ^ ((~A[4][2][8]) & A[0][2][8]);
   assign A_chi[2][3][9]     = A[3][2][9] ^ ((~A[4][2][9]) & A[0][2][9]);
   assign A_chi[2][3][10]     = A[3][2][10] ^ ((~A[4][2][10]) & A[0][2][10]);
   assign A_chi[2][3][11]     = A[3][2][11] ^ ((~A[4][2][11]) & A[0][2][11]);
   assign A_chi[2][3][12]     = A[3][2][12] ^ ((~A[4][2][12]) & A[0][2][12]);
   assign A_chi[2][3][13]     = A[3][2][13] ^ ((~A[4][2][13]) & A[0][2][13]);
   assign A_chi[2][3][14]     = A[3][2][14] ^ ((~A[4][2][14]) & A[0][2][14]);
   assign A_chi[2][3][15]     = A[3][2][15] ^ ((~A[4][2][15]) & A[0][2][15]);
   assign A_chi[2][3][16]     = A[3][2][16] ^ ((~A[4][2][16]) & A[0][2][16]);
   assign A_chi[2][3][17]     = A[3][2][17] ^ ((~A[4][2][17]) & A[0][2][17]);
   assign A_chi[2][3][18]     = A[3][2][18] ^ ((~A[4][2][18]) & A[0][2][18]);
   assign A_chi[2][3][19]     = A[3][2][19] ^ ((~A[4][2][19]) & A[0][2][19]);
   assign A_chi[2][3][20]     = A[3][2][20] ^ ((~A[4][2][20]) & A[0][2][20]);
   assign A_chi[2][3][21]     = A[3][2][21] ^ ((~A[4][2][21]) & A[0][2][21]);
   assign A_chi[2][3][22]     = A[3][2][22] ^ ((~A[4][2][22]) & A[0][2][22]);
   assign A_chi[2][3][23]     = A[3][2][23] ^ ((~A[4][2][23]) & A[0][2][23]);
   assign A_chi[2][3][24]     = A[3][2][24] ^ ((~A[4][2][24]) & A[0][2][24]);
   assign A_chi[2][3][25]     = A[3][2][25] ^ ((~A[4][2][25]) & A[0][2][25]);
   assign A_chi[2][3][26]     = A[3][2][26] ^ ((~A[4][2][26]) & A[0][2][26]);
   assign A_chi[2][3][27]     = A[3][2][27] ^ ((~A[4][2][27]) & A[0][2][27]);
   assign A_chi[2][3][28]     = A[3][2][28] ^ ((~A[4][2][28]) & A[0][2][28]);
   assign A_chi[2][3][29]     = A[3][2][29] ^ ((~A[4][2][29]) & A[0][2][29]);
   assign A_chi[2][3][30]     = A[3][2][30] ^ ((~A[4][2][30]) & A[0][2][30]);
   assign A_chi[2][3][31]     = A[3][2][31] ^ ((~A[4][2][31]) & A[0][2][31]);
   assign A_chi[2][3][32]     = A[3][2][32] ^ ((~A[4][2][32]) & A[0][2][32]);
   assign A_chi[2][3][33]     = A[3][2][33] ^ ((~A[4][2][33]) & A[0][2][33]);
   assign A_chi[2][3][34]     = A[3][2][34] ^ ((~A[4][2][34]) & A[0][2][34]);
   assign A_chi[2][3][35]     = A[3][2][35] ^ ((~A[4][2][35]) & A[0][2][35]);
   assign A_chi[2][3][36]     = A[3][2][36] ^ ((~A[4][2][36]) & A[0][2][36]);
   assign A_chi[2][3][37]     = A[3][2][37] ^ ((~A[4][2][37]) & A[0][2][37]);
   assign A_chi[2][3][38]     = A[3][2][38] ^ ((~A[4][2][38]) & A[0][2][38]);
   assign A_chi[2][3][39]     = A[3][2][39] ^ ((~A[4][2][39]) & A[0][2][39]);
   assign A_chi[2][3][40]     = A[3][2][40] ^ ((~A[4][2][40]) & A[0][2][40]);
   assign A_chi[2][3][41]     = A[3][2][41] ^ ((~A[4][2][41]) & A[0][2][41]);
   assign A_chi[2][3][42]     = A[3][2][42] ^ ((~A[4][2][42]) & A[0][2][42]);
   assign A_chi[2][3][43]     = A[3][2][43] ^ ((~A[4][2][43]) & A[0][2][43]);
   assign A_chi[2][3][44]     = A[3][2][44] ^ ((~A[4][2][44]) & A[0][2][44]);
   assign A_chi[2][3][45]     = A[3][2][45] ^ ((~A[4][2][45]) & A[0][2][45]);
   assign A_chi[2][3][46]     = A[3][2][46] ^ ((~A[4][2][46]) & A[0][2][46]);
   assign A_chi[2][3][47]     = A[3][2][47] ^ ((~A[4][2][47]) & A[0][2][47]);
   assign A_chi[2][3][48]     = A[3][2][48] ^ ((~A[4][2][48]) & A[0][2][48]);
   assign A_chi[2][3][49]     = A[3][2][49] ^ ((~A[4][2][49]) & A[0][2][49]);
   assign A_chi[2][3][50]     = A[3][2][50] ^ ((~A[4][2][50]) & A[0][2][50]);
   assign A_chi[2][3][51]     = A[3][2][51] ^ ((~A[4][2][51]) & A[0][2][51]);
   assign A_chi[2][3][52]     = A[3][2][52] ^ ((~A[4][2][52]) & A[0][2][52]);
   assign A_chi[2][3][53]     = A[3][2][53] ^ ((~A[4][2][53]) & A[0][2][53]);
   assign A_chi[2][3][54]     = A[3][2][54] ^ ((~A[4][2][54]) & A[0][2][54]);
   assign A_chi[2][3][55]     = A[3][2][55] ^ ((~A[4][2][55]) & A[0][2][55]);
   assign A_chi[2][3][56]     = A[3][2][56] ^ ((~A[4][2][56]) & A[0][2][56]);
   assign A_chi[2][3][57]     = A[3][2][57] ^ ((~A[4][2][57]) & A[0][2][57]);
   assign A_chi[2][3][58]     = A[3][2][58] ^ ((~A[4][2][58]) & A[0][2][58]);
   assign A_chi[2][3][59]     = A[3][2][59] ^ ((~A[4][2][59]) & A[0][2][59]);
   assign A_chi[2][3][60]     = A[3][2][60] ^ ((~A[4][2][60]) & A[0][2][60]);
   assign A_chi[2][3][61]     = A[3][2][61] ^ ((~A[4][2][61]) & A[0][2][61]);
   assign A_chi[2][3][62]     = A[3][2][62] ^ ((~A[4][2][62]) & A[0][2][62]);
   assign A_chi[2][3][63]     = A[3][2][63] ^ ((~A[4][2][63]) & A[0][2][63]);
   assign A_chi[2][4][0]     = A[4][2][0] ^ ((~A[0][2][0]) & A[1][2][0]);
   assign A_chi[2][4][1]     = A[4][2][1] ^ ((~A[0][2][1]) & A[1][2][1]);
   assign A_chi[2][4][2]     = A[4][2][2] ^ ((~A[0][2][2]) & A[1][2][2]);
   assign A_chi[2][4][3]     = A[4][2][3] ^ ((~A[0][2][3]) & A[1][2][3]);
   assign A_chi[2][4][4]     = A[4][2][4] ^ ((~A[0][2][4]) & A[1][2][4]);
   assign A_chi[2][4][5]     = A[4][2][5] ^ ((~A[0][2][5]) & A[1][2][5]);
   assign A_chi[2][4][6]     = A[4][2][6] ^ ((~A[0][2][6]) & A[1][2][6]);
   assign A_chi[2][4][7]     = A[4][2][7] ^ ((~A[0][2][7]) & A[1][2][7]);
   assign A_chi[2][4][8]     = A[4][2][8] ^ ((~A[0][2][8]) & A[1][2][8]);
   assign A_chi[2][4][9]     = A[4][2][9] ^ ((~A[0][2][9]) & A[1][2][9]);
   assign A_chi[2][4][10]     = A[4][2][10] ^ ((~A[0][2][10]) & A[1][2][10]);
   assign A_chi[2][4][11]     = A[4][2][11] ^ ((~A[0][2][11]) & A[1][2][11]);
   assign A_chi[2][4][12]     = A[4][2][12] ^ ((~A[0][2][12]) & A[1][2][12]);
   assign A_chi[2][4][13]     = A[4][2][13] ^ ((~A[0][2][13]) & A[1][2][13]);
   assign A_chi[2][4][14]     = A[4][2][14] ^ ((~A[0][2][14]) & A[1][2][14]);
   assign A_chi[2][4][15]     = A[4][2][15] ^ ((~A[0][2][15]) & A[1][2][15]);
   assign A_chi[2][4][16]     = A[4][2][16] ^ ((~A[0][2][16]) & A[1][2][16]);
   assign A_chi[2][4][17]     = A[4][2][17] ^ ((~A[0][2][17]) & A[1][2][17]);
   assign A_chi[2][4][18]     = A[4][2][18] ^ ((~A[0][2][18]) & A[1][2][18]);
   assign A_chi[2][4][19]     = A[4][2][19] ^ ((~A[0][2][19]) & A[1][2][19]);
   assign A_chi[2][4][20]     = A[4][2][20] ^ ((~A[0][2][20]) & A[1][2][20]);
   assign A_chi[2][4][21]     = A[4][2][21] ^ ((~A[0][2][21]) & A[1][2][21]);
   assign A_chi[2][4][22]     = A[4][2][22] ^ ((~A[0][2][22]) & A[1][2][22]);
   assign A_chi[2][4][23]     = A[4][2][23] ^ ((~A[0][2][23]) & A[1][2][23]);
   assign A_chi[2][4][24]     = A[4][2][24] ^ ((~A[0][2][24]) & A[1][2][24]);
   assign A_chi[2][4][25]     = A[4][2][25] ^ ((~A[0][2][25]) & A[1][2][25]);
   assign A_chi[2][4][26]     = A[4][2][26] ^ ((~A[0][2][26]) & A[1][2][26]);
   assign A_chi[2][4][27]     = A[4][2][27] ^ ((~A[0][2][27]) & A[1][2][27]);
   assign A_chi[2][4][28]     = A[4][2][28] ^ ((~A[0][2][28]) & A[1][2][28]);
   assign A_chi[2][4][29]     = A[4][2][29] ^ ((~A[0][2][29]) & A[1][2][29]);
   assign A_chi[2][4][30]     = A[4][2][30] ^ ((~A[0][2][30]) & A[1][2][30]);
   assign A_chi[2][4][31]     = A[4][2][31] ^ ((~A[0][2][31]) & A[1][2][31]);
   assign A_chi[2][4][32]     = A[4][2][32] ^ ((~A[0][2][32]) & A[1][2][32]);
   assign A_chi[2][4][33]     = A[4][2][33] ^ ((~A[0][2][33]) & A[1][2][33]);
   assign A_chi[2][4][34]     = A[4][2][34] ^ ((~A[0][2][34]) & A[1][2][34]);
   assign A_chi[2][4][35]     = A[4][2][35] ^ ((~A[0][2][35]) & A[1][2][35]);
   assign A_chi[2][4][36]     = A[4][2][36] ^ ((~A[0][2][36]) & A[1][2][36]);
   assign A_chi[2][4][37]     = A[4][2][37] ^ ((~A[0][2][37]) & A[1][2][37]);
   assign A_chi[2][4][38]     = A[4][2][38] ^ ((~A[0][2][38]) & A[1][2][38]);
   assign A_chi[2][4][39]     = A[4][2][39] ^ ((~A[0][2][39]) & A[1][2][39]);
   assign A_chi[2][4][40]     = A[4][2][40] ^ ((~A[0][2][40]) & A[1][2][40]);
   assign A_chi[2][4][41]     = A[4][2][41] ^ ((~A[0][2][41]) & A[1][2][41]);
   assign A_chi[2][4][42]     = A[4][2][42] ^ ((~A[0][2][42]) & A[1][2][42]);
   assign A_chi[2][4][43]     = A[4][2][43] ^ ((~A[0][2][43]) & A[1][2][43]);
   assign A_chi[2][4][44]     = A[4][2][44] ^ ((~A[0][2][44]) & A[1][2][44]);
   assign A_chi[2][4][45]     = A[4][2][45] ^ ((~A[0][2][45]) & A[1][2][45]);
   assign A_chi[2][4][46]     = A[4][2][46] ^ ((~A[0][2][46]) & A[1][2][46]);
   assign A_chi[2][4][47]     = A[4][2][47] ^ ((~A[0][2][47]) & A[1][2][47]);
   assign A_chi[2][4][48]     = A[4][2][48] ^ ((~A[0][2][48]) & A[1][2][48]);
   assign A_chi[2][4][49]     = A[4][2][49] ^ ((~A[0][2][49]) & A[1][2][49]);
   assign A_chi[2][4][50]     = A[4][2][50] ^ ((~A[0][2][50]) & A[1][2][50]);
   assign A_chi[2][4][51]     = A[4][2][51] ^ ((~A[0][2][51]) & A[1][2][51]);
   assign A_chi[2][4][52]     = A[4][2][52] ^ ((~A[0][2][52]) & A[1][2][52]);
   assign A_chi[2][4][53]     = A[4][2][53] ^ ((~A[0][2][53]) & A[1][2][53]);
   assign A_chi[2][4][54]     = A[4][2][54] ^ ((~A[0][2][54]) & A[1][2][54]);
   assign A_chi[2][4][55]     = A[4][2][55] ^ ((~A[0][2][55]) & A[1][2][55]);
   assign A_chi[2][4][56]     = A[4][2][56] ^ ((~A[0][2][56]) & A[1][2][56]);
   assign A_chi[2][4][57]     = A[4][2][57] ^ ((~A[0][2][57]) & A[1][2][57]);
   assign A_chi[2][4][58]     = A[4][2][58] ^ ((~A[0][2][58]) & A[1][2][58]);
   assign A_chi[2][4][59]     = A[4][2][59] ^ ((~A[0][2][59]) & A[1][2][59]);
   assign A_chi[2][4][60]     = A[4][2][60] ^ ((~A[0][2][60]) & A[1][2][60]);
   assign A_chi[2][4][61]     = A[4][2][61] ^ ((~A[0][2][61]) & A[1][2][61]);
   assign A_chi[2][4][62]     = A[4][2][62] ^ ((~A[0][2][62]) & A[1][2][62]);
   assign A_chi[2][4][63]     = A[4][2][63] ^ ((~A[0][2][63]) & A[1][2][63]);
   assign A_chi[3][0][0]     = A[0][3][0] ^ ((~A[1][3][0]) & A[2][3][0]);
   assign A_chi[3][0][1]     = A[0][3][1] ^ ((~A[1][3][1]) & A[2][3][1]);
   assign A_chi[3][0][2]     = A[0][3][2] ^ ((~A[1][3][2]) & A[2][3][2]);
   assign A_chi[3][0][3]     = A[0][3][3] ^ ((~A[1][3][3]) & A[2][3][3]);
   assign A_chi[3][0][4]     = A[0][3][4] ^ ((~A[1][3][4]) & A[2][3][4]);
   assign A_chi[3][0][5]     = A[0][3][5] ^ ((~A[1][3][5]) & A[2][3][5]);
   assign A_chi[3][0][6]     = A[0][3][6] ^ ((~A[1][3][6]) & A[2][3][6]);
   assign A_chi[3][0][7]     = A[0][3][7] ^ ((~A[1][3][7]) & A[2][3][7]);
   assign A_chi[3][0][8]     = A[0][3][8] ^ ((~A[1][3][8]) & A[2][3][8]);
   assign A_chi[3][0][9]     = A[0][3][9] ^ ((~A[1][3][9]) & A[2][3][9]);
   assign A_chi[3][0][10]     = A[0][3][10] ^ ((~A[1][3][10]) & A[2][3][10]);
   assign A_chi[3][0][11]     = A[0][3][11] ^ ((~A[1][3][11]) & A[2][3][11]);
   assign A_chi[3][0][12]     = A[0][3][12] ^ ((~A[1][3][12]) & A[2][3][12]);
   assign A_chi[3][0][13]     = A[0][3][13] ^ ((~A[1][3][13]) & A[2][3][13]);
   assign A_chi[3][0][14]     = A[0][3][14] ^ ((~A[1][3][14]) & A[2][3][14]);
   assign A_chi[3][0][15]     = A[0][3][15] ^ ((~A[1][3][15]) & A[2][3][15]);
   assign A_chi[3][0][16]     = A[0][3][16] ^ ((~A[1][3][16]) & A[2][3][16]);
   assign A_chi[3][0][17]     = A[0][3][17] ^ ((~A[1][3][17]) & A[2][3][17]);
   assign A_chi[3][0][18]     = A[0][3][18] ^ ((~A[1][3][18]) & A[2][3][18]);
   assign A_chi[3][0][19]     = A[0][3][19] ^ ((~A[1][3][19]) & A[2][3][19]);
   assign A_chi[3][0][20]     = A[0][3][20] ^ ((~A[1][3][20]) & A[2][3][20]);
   assign A_chi[3][0][21]     = A[0][3][21] ^ ((~A[1][3][21]) & A[2][3][21]);
   assign A_chi[3][0][22]     = A[0][3][22] ^ ((~A[1][3][22]) & A[2][3][22]);
   assign A_chi[3][0][23]     = A[0][3][23] ^ ((~A[1][3][23]) & A[2][3][23]);
   assign A_chi[3][0][24]     = A[0][3][24] ^ ((~A[1][3][24]) & A[2][3][24]);
   assign A_chi[3][0][25]     = A[0][3][25] ^ ((~A[1][3][25]) & A[2][3][25]);
   assign A_chi[3][0][26]     = A[0][3][26] ^ ((~A[1][3][26]) & A[2][3][26]);
   assign A_chi[3][0][27]     = A[0][3][27] ^ ((~A[1][3][27]) & A[2][3][27]);
   assign A_chi[3][0][28]     = A[0][3][28] ^ ((~A[1][3][28]) & A[2][3][28]);
   assign A_chi[3][0][29]     = A[0][3][29] ^ ((~A[1][3][29]) & A[2][3][29]);
   assign A_chi[3][0][30]     = A[0][3][30] ^ ((~A[1][3][30]) & A[2][3][30]);
   assign A_chi[3][0][31]     = A[0][3][31] ^ ((~A[1][3][31]) & A[2][3][31]);
   assign A_chi[3][0][32]     = A[0][3][32] ^ ((~A[1][3][32]) & A[2][3][32]);
   assign A_chi[3][0][33]     = A[0][3][33] ^ ((~A[1][3][33]) & A[2][3][33]);
   assign A_chi[3][0][34]     = A[0][3][34] ^ ((~A[1][3][34]) & A[2][3][34]);
   assign A_chi[3][0][35]     = A[0][3][35] ^ ((~A[1][3][35]) & A[2][3][35]);
   assign A_chi[3][0][36]     = A[0][3][36] ^ ((~A[1][3][36]) & A[2][3][36]);
   assign A_chi[3][0][37]     = A[0][3][37] ^ ((~A[1][3][37]) & A[2][3][37]);
   assign A_chi[3][0][38]     = A[0][3][38] ^ ((~A[1][3][38]) & A[2][3][38]);
   assign A_chi[3][0][39]     = A[0][3][39] ^ ((~A[1][3][39]) & A[2][3][39]);
   assign A_chi[3][0][40]     = A[0][3][40] ^ ((~A[1][3][40]) & A[2][3][40]);
   assign A_chi[3][0][41]     = A[0][3][41] ^ ((~A[1][3][41]) & A[2][3][41]);
   assign A_chi[3][0][42]     = A[0][3][42] ^ ((~A[1][3][42]) & A[2][3][42]);
   assign A_chi[3][0][43]     = A[0][3][43] ^ ((~A[1][3][43]) & A[2][3][43]);
   assign A_chi[3][0][44]     = A[0][3][44] ^ ((~A[1][3][44]) & A[2][3][44]);
   assign A_chi[3][0][45]     = A[0][3][45] ^ ((~A[1][3][45]) & A[2][3][45]);
   assign A_chi[3][0][46]     = A[0][3][46] ^ ((~A[1][3][46]) & A[2][3][46]);
   assign A_chi[3][0][47]     = A[0][3][47] ^ ((~A[1][3][47]) & A[2][3][47]);
   assign A_chi[3][0][48]     = A[0][3][48] ^ ((~A[1][3][48]) & A[2][3][48]);
   assign A_chi[3][0][49]     = A[0][3][49] ^ ((~A[1][3][49]) & A[2][3][49]);
   assign A_chi[3][0][50]     = A[0][3][50] ^ ((~A[1][3][50]) & A[2][3][50]);
   assign A_chi[3][0][51]     = A[0][3][51] ^ ((~A[1][3][51]) & A[2][3][51]);
   assign A_chi[3][0][52]     = A[0][3][52] ^ ((~A[1][3][52]) & A[2][3][52]);
   assign A_chi[3][0][53]     = A[0][3][53] ^ ((~A[1][3][53]) & A[2][3][53]);
   assign A_chi[3][0][54]     = A[0][3][54] ^ ((~A[1][3][54]) & A[2][3][54]);
   assign A_chi[3][0][55]     = A[0][3][55] ^ ((~A[1][3][55]) & A[2][3][55]);
   assign A_chi[3][0][56]     = A[0][3][56] ^ ((~A[1][3][56]) & A[2][3][56]);
   assign A_chi[3][0][57]     = A[0][3][57] ^ ((~A[1][3][57]) & A[2][3][57]);
   assign A_chi[3][0][58]     = A[0][3][58] ^ ((~A[1][3][58]) & A[2][3][58]);
   assign A_chi[3][0][59]     = A[0][3][59] ^ ((~A[1][3][59]) & A[2][3][59]);
   assign A_chi[3][0][60]     = A[0][3][60] ^ ((~A[1][3][60]) & A[2][3][60]);
   assign A_chi[3][0][61]     = A[0][3][61] ^ ((~A[1][3][61]) & A[2][3][61]);
   assign A_chi[3][0][62]     = A[0][3][62] ^ ((~A[1][3][62]) & A[2][3][62]);
   assign A_chi[3][0][63]     = A[0][3][63] ^ ((~A[1][3][63]) & A[2][3][63]);
   assign A_chi[3][1][0]     = A[1][3][0] ^ ((~A[2][3][0]) & A[3][3][0]);
   assign A_chi[3][1][1]     = A[1][3][1] ^ ((~A[2][3][1]) & A[3][3][1]);
   assign A_chi[3][1][2]     = A[1][3][2] ^ ((~A[2][3][2]) & A[3][3][2]);
   assign A_chi[3][1][3]     = A[1][3][3] ^ ((~A[2][3][3]) & A[3][3][3]);
   assign A_chi[3][1][4]     = A[1][3][4] ^ ((~A[2][3][4]) & A[3][3][4]);
   assign A_chi[3][1][5]     = A[1][3][5] ^ ((~A[2][3][5]) & A[3][3][5]);
   assign A_chi[3][1][6]     = A[1][3][6] ^ ((~A[2][3][6]) & A[3][3][6]);
   assign A_chi[3][1][7]     = A[1][3][7] ^ ((~A[2][3][7]) & A[3][3][7]);
   assign A_chi[3][1][8]     = A[1][3][8] ^ ((~A[2][3][8]) & A[3][3][8]);
   assign A_chi[3][1][9]     = A[1][3][9] ^ ((~A[2][3][9]) & A[3][3][9]);
   assign A_chi[3][1][10]     = A[1][3][10] ^ ((~A[2][3][10]) & A[3][3][10]);
   assign A_chi[3][1][11]     = A[1][3][11] ^ ((~A[2][3][11]) & A[3][3][11]);
   assign A_chi[3][1][12]     = A[1][3][12] ^ ((~A[2][3][12]) & A[3][3][12]);
   assign A_chi[3][1][13]     = A[1][3][13] ^ ((~A[2][3][13]) & A[3][3][13]);
   assign A_chi[3][1][14]     = A[1][3][14] ^ ((~A[2][3][14]) & A[3][3][14]);
   assign A_chi[3][1][15]     = A[1][3][15] ^ ((~A[2][3][15]) & A[3][3][15]);
   assign A_chi[3][1][16]     = A[1][3][16] ^ ((~A[2][3][16]) & A[3][3][16]);
   assign A_chi[3][1][17]     = A[1][3][17] ^ ((~A[2][3][17]) & A[3][3][17]);
   assign A_chi[3][1][18]     = A[1][3][18] ^ ((~A[2][3][18]) & A[3][3][18]);
   assign A_chi[3][1][19]     = A[1][3][19] ^ ((~A[2][3][19]) & A[3][3][19]);
   assign A_chi[3][1][20]     = A[1][3][20] ^ ((~A[2][3][20]) & A[3][3][20]);
   assign A_chi[3][1][21]     = A[1][3][21] ^ ((~A[2][3][21]) & A[3][3][21]);
   assign A_chi[3][1][22]     = A[1][3][22] ^ ((~A[2][3][22]) & A[3][3][22]);
   assign A_chi[3][1][23]     = A[1][3][23] ^ ((~A[2][3][23]) & A[3][3][23]);
   assign A_chi[3][1][24]     = A[1][3][24] ^ ((~A[2][3][24]) & A[3][3][24]);
   assign A_chi[3][1][25]     = A[1][3][25] ^ ((~A[2][3][25]) & A[3][3][25]);
   assign A_chi[3][1][26]     = A[1][3][26] ^ ((~A[2][3][26]) & A[3][3][26]);
   assign A_chi[3][1][27]     = A[1][3][27] ^ ((~A[2][3][27]) & A[3][3][27]);
   assign A_chi[3][1][28]     = A[1][3][28] ^ ((~A[2][3][28]) & A[3][3][28]);
   assign A_chi[3][1][29]     = A[1][3][29] ^ ((~A[2][3][29]) & A[3][3][29]);
   assign A_chi[3][1][30]     = A[1][3][30] ^ ((~A[2][3][30]) & A[3][3][30]);
   assign A_chi[3][1][31]     = A[1][3][31] ^ ((~A[2][3][31]) & A[3][3][31]);
   assign A_chi[3][1][32]     = A[1][3][32] ^ ((~A[2][3][32]) & A[3][3][32]);
   assign A_chi[3][1][33]     = A[1][3][33] ^ ((~A[2][3][33]) & A[3][3][33]);
   assign A_chi[3][1][34]     = A[1][3][34] ^ ((~A[2][3][34]) & A[3][3][34]);
   assign A_chi[3][1][35]     = A[1][3][35] ^ ((~A[2][3][35]) & A[3][3][35]);
   assign A_chi[3][1][36]     = A[1][3][36] ^ ((~A[2][3][36]) & A[3][3][36]);
   assign A_chi[3][1][37]     = A[1][3][37] ^ ((~A[2][3][37]) & A[3][3][37]);
   assign A_chi[3][1][38]     = A[1][3][38] ^ ((~A[2][3][38]) & A[3][3][38]);
   assign A_chi[3][1][39]     = A[1][3][39] ^ ((~A[2][3][39]) & A[3][3][39]);
   assign A_chi[3][1][40]     = A[1][3][40] ^ ((~A[2][3][40]) & A[3][3][40]);
   assign A_chi[3][1][41]     = A[1][3][41] ^ ((~A[2][3][41]) & A[3][3][41]);
   assign A_chi[3][1][42]     = A[1][3][42] ^ ((~A[2][3][42]) & A[3][3][42]);
   assign A_chi[3][1][43]     = A[1][3][43] ^ ((~A[2][3][43]) & A[3][3][43]);
   assign A_chi[3][1][44]     = A[1][3][44] ^ ((~A[2][3][44]) & A[3][3][44]);
   assign A_chi[3][1][45]     = A[1][3][45] ^ ((~A[2][3][45]) & A[3][3][45]);
   assign A_chi[3][1][46]     = A[1][3][46] ^ ((~A[2][3][46]) & A[3][3][46]);
   assign A_chi[3][1][47]     = A[1][3][47] ^ ((~A[2][3][47]) & A[3][3][47]);
   assign A_chi[3][1][48]     = A[1][3][48] ^ ((~A[2][3][48]) & A[3][3][48]);
   assign A_chi[3][1][49]     = A[1][3][49] ^ ((~A[2][3][49]) & A[3][3][49]);
   assign A_chi[3][1][50]     = A[1][3][50] ^ ((~A[2][3][50]) & A[3][3][50]);
   assign A_chi[3][1][51]     = A[1][3][51] ^ ((~A[2][3][51]) & A[3][3][51]);
   assign A_chi[3][1][52]     = A[1][3][52] ^ ((~A[2][3][52]) & A[3][3][52]);
   assign A_chi[3][1][53]     = A[1][3][53] ^ ((~A[2][3][53]) & A[3][3][53]);
   assign A_chi[3][1][54]     = A[1][3][54] ^ ((~A[2][3][54]) & A[3][3][54]);
   assign A_chi[3][1][55]     = A[1][3][55] ^ ((~A[2][3][55]) & A[3][3][55]);
   assign A_chi[3][1][56]     = A[1][3][56] ^ ((~A[2][3][56]) & A[3][3][56]);
   assign A_chi[3][1][57]     = A[1][3][57] ^ ((~A[2][3][57]) & A[3][3][57]);
   assign A_chi[3][1][58]     = A[1][3][58] ^ ((~A[2][3][58]) & A[3][3][58]);
   assign A_chi[3][1][59]     = A[1][3][59] ^ ((~A[2][3][59]) & A[3][3][59]);
   assign A_chi[3][1][60]     = A[1][3][60] ^ ((~A[2][3][60]) & A[3][3][60]);
   assign A_chi[3][1][61]     = A[1][3][61] ^ ((~A[2][3][61]) & A[3][3][61]);
   assign A_chi[3][1][62]     = A[1][3][62] ^ ((~A[2][3][62]) & A[3][3][62]);
   assign A_chi[3][1][63]     = A[1][3][63] ^ ((~A[2][3][63]) & A[3][3][63]);
   assign A_chi[3][2][0]     = A[2][3][0] ^ ((~A[3][3][0]) & A[4][3][0]);
   assign A_chi[3][2][1]     = A[2][3][1] ^ ((~A[3][3][1]) & A[4][3][1]);
   assign A_chi[3][2][2]     = A[2][3][2] ^ ((~A[3][3][2]) & A[4][3][2]);
   assign A_chi[3][2][3]     = A[2][3][3] ^ ((~A[3][3][3]) & A[4][3][3]);
   assign A_chi[3][2][4]     = A[2][3][4] ^ ((~A[3][3][4]) & A[4][3][4]);
   assign A_chi[3][2][5]     = A[2][3][5] ^ ((~A[3][3][5]) & A[4][3][5]);
   assign A_chi[3][2][6]     = A[2][3][6] ^ ((~A[3][3][6]) & A[4][3][6]);
   assign A_chi[3][2][7]     = A[2][3][7] ^ ((~A[3][3][7]) & A[4][3][7]);
   assign A_chi[3][2][8]     = A[2][3][8] ^ ((~A[3][3][8]) & A[4][3][8]);
   assign A_chi[3][2][9]     = A[2][3][9] ^ ((~A[3][3][9]) & A[4][3][9]);
   assign A_chi[3][2][10]     = A[2][3][10] ^ ((~A[3][3][10]) & A[4][3][10]);
   assign A_chi[3][2][11]     = A[2][3][11] ^ ((~A[3][3][11]) & A[4][3][11]);
   assign A_chi[3][2][12]     = A[2][3][12] ^ ((~A[3][3][12]) & A[4][3][12]);
   assign A_chi[3][2][13]     = A[2][3][13] ^ ((~A[3][3][13]) & A[4][3][13]);
   assign A_chi[3][2][14]     = A[2][3][14] ^ ((~A[3][3][14]) & A[4][3][14]);
   assign A_chi[3][2][15]     = A[2][3][15] ^ ((~A[3][3][15]) & A[4][3][15]);
   assign A_chi[3][2][16]     = A[2][3][16] ^ ((~A[3][3][16]) & A[4][3][16]);
   assign A_chi[3][2][17]     = A[2][3][17] ^ ((~A[3][3][17]) & A[4][3][17]);
   assign A_chi[3][2][18]     = A[2][3][18] ^ ((~A[3][3][18]) & A[4][3][18]);
   assign A_chi[3][2][19]     = A[2][3][19] ^ ((~A[3][3][19]) & A[4][3][19]);
   assign A_chi[3][2][20]     = A[2][3][20] ^ ((~A[3][3][20]) & A[4][3][20]);
   assign A_chi[3][2][21]     = A[2][3][21] ^ ((~A[3][3][21]) & A[4][3][21]);
   assign A_chi[3][2][22]     = A[2][3][22] ^ ((~A[3][3][22]) & A[4][3][22]);
   assign A_chi[3][2][23]     = A[2][3][23] ^ ((~A[3][3][23]) & A[4][3][23]);
   assign A_chi[3][2][24]     = A[2][3][24] ^ ((~A[3][3][24]) & A[4][3][24]);
   assign A_chi[3][2][25]     = A[2][3][25] ^ ((~A[3][3][25]) & A[4][3][25]);
   assign A_chi[3][2][26]     = A[2][3][26] ^ ((~A[3][3][26]) & A[4][3][26]);
   assign A_chi[3][2][27]     = A[2][3][27] ^ ((~A[3][3][27]) & A[4][3][27]);
   assign A_chi[3][2][28]     = A[2][3][28] ^ ((~A[3][3][28]) & A[4][3][28]);
   assign A_chi[3][2][29]     = A[2][3][29] ^ ((~A[3][3][29]) & A[4][3][29]);
   assign A_chi[3][2][30]     = A[2][3][30] ^ ((~A[3][3][30]) & A[4][3][30]);
   assign A_chi[3][2][31]     = A[2][3][31] ^ ((~A[3][3][31]) & A[4][3][31]);
   assign A_chi[3][2][32]     = A[2][3][32] ^ ((~A[3][3][32]) & A[4][3][32]);
   assign A_chi[3][2][33]     = A[2][3][33] ^ ((~A[3][3][33]) & A[4][3][33]);
   assign A_chi[3][2][34]     = A[2][3][34] ^ ((~A[3][3][34]) & A[4][3][34]);
   assign A_chi[3][2][35]     = A[2][3][35] ^ ((~A[3][3][35]) & A[4][3][35]);
   assign A_chi[3][2][36]     = A[2][3][36] ^ ((~A[3][3][36]) & A[4][3][36]);
   assign A_chi[3][2][37]     = A[2][3][37] ^ ((~A[3][3][37]) & A[4][3][37]);
   assign A_chi[3][2][38]     = A[2][3][38] ^ ((~A[3][3][38]) & A[4][3][38]);
   assign A_chi[3][2][39]     = A[2][3][39] ^ ((~A[3][3][39]) & A[4][3][39]);
   assign A_chi[3][2][40]     = A[2][3][40] ^ ((~A[3][3][40]) & A[4][3][40]);
   assign A_chi[3][2][41]     = A[2][3][41] ^ ((~A[3][3][41]) & A[4][3][41]);
   assign A_chi[3][2][42]     = A[2][3][42] ^ ((~A[3][3][42]) & A[4][3][42]);
   assign A_chi[3][2][43]     = A[2][3][43] ^ ((~A[3][3][43]) & A[4][3][43]);
   assign A_chi[3][2][44]     = A[2][3][44] ^ ((~A[3][3][44]) & A[4][3][44]);
   assign A_chi[3][2][45]     = A[2][3][45] ^ ((~A[3][3][45]) & A[4][3][45]);
   assign A_chi[3][2][46]     = A[2][3][46] ^ ((~A[3][3][46]) & A[4][3][46]);
   assign A_chi[3][2][47]     = A[2][3][47] ^ ((~A[3][3][47]) & A[4][3][47]);
   assign A_chi[3][2][48]     = A[2][3][48] ^ ((~A[3][3][48]) & A[4][3][48]);
   assign A_chi[3][2][49]     = A[2][3][49] ^ ((~A[3][3][49]) & A[4][3][49]);
   assign A_chi[3][2][50]     = A[2][3][50] ^ ((~A[3][3][50]) & A[4][3][50]);
   assign A_chi[3][2][51]     = A[2][3][51] ^ ((~A[3][3][51]) & A[4][3][51]);
   assign A_chi[3][2][52]     = A[2][3][52] ^ ((~A[3][3][52]) & A[4][3][52]);
   assign A_chi[3][2][53]     = A[2][3][53] ^ ((~A[3][3][53]) & A[4][3][53]);
   assign A_chi[3][2][54]     = A[2][3][54] ^ ((~A[3][3][54]) & A[4][3][54]);
   assign A_chi[3][2][55]     = A[2][3][55] ^ ((~A[3][3][55]) & A[4][3][55]);
   assign A_chi[3][2][56]     = A[2][3][56] ^ ((~A[3][3][56]) & A[4][3][56]);
   assign A_chi[3][2][57]     = A[2][3][57] ^ ((~A[3][3][57]) & A[4][3][57]);
   assign A_chi[3][2][58]     = A[2][3][58] ^ ((~A[3][3][58]) & A[4][3][58]);
   assign A_chi[3][2][59]     = A[2][3][59] ^ ((~A[3][3][59]) & A[4][3][59]);
   assign A_chi[3][2][60]     = A[2][3][60] ^ ((~A[3][3][60]) & A[4][3][60]);
   assign A_chi[3][2][61]     = A[2][3][61] ^ ((~A[3][3][61]) & A[4][3][61]);
   assign A_chi[3][2][62]     = A[2][3][62] ^ ((~A[3][3][62]) & A[4][3][62]);
   assign A_chi[3][2][63]     = A[2][3][63] ^ ((~A[3][3][63]) & A[4][3][63]);
   assign A_chi[3][3][0]     = A[3][3][0] ^ ((~A[4][3][0]) & A[0][3][0]);
   assign A_chi[3][3][1]     = A[3][3][1] ^ ((~A[4][3][1]) & A[0][3][1]);
   assign A_chi[3][3][2]     = A[3][3][2] ^ ((~A[4][3][2]) & A[0][3][2]);
   assign A_chi[3][3][3]     = A[3][3][3] ^ ((~A[4][3][3]) & A[0][3][3]);
   assign A_chi[3][3][4]     = A[3][3][4] ^ ((~A[4][3][4]) & A[0][3][4]);
   assign A_chi[3][3][5]     = A[3][3][5] ^ ((~A[4][3][5]) & A[0][3][5]);
   assign A_chi[3][3][6]     = A[3][3][6] ^ ((~A[4][3][6]) & A[0][3][6]);
   assign A_chi[3][3][7]     = A[3][3][7] ^ ((~A[4][3][7]) & A[0][3][7]);
   assign A_chi[3][3][8]     = A[3][3][8] ^ ((~A[4][3][8]) & A[0][3][8]);
   assign A_chi[3][3][9]     = A[3][3][9] ^ ((~A[4][3][9]) & A[0][3][9]);
   assign A_chi[3][3][10]     = A[3][3][10] ^ ((~A[4][3][10]) & A[0][3][10]);
   assign A_chi[3][3][11]     = A[3][3][11] ^ ((~A[4][3][11]) & A[0][3][11]);
   assign A_chi[3][3][12]     = A[3][3][12] ^ ((~A[4][3][12]) & A[0][3][12]);
   assign A_chi[3][3][13]     = A[3][3][13] ^ ((~A[4][3][13]) & A[0][3][13]);
   assign A_chi[3][3][14]     = A[3][3][14] ^ ((~A[4][3][14]) & A[0][3][14]);
   assign A_chi[3][3][15]     = A[3][3][15] ^ ((~A[4][3][15]) & A[0][3][15]);
   assign A_chi[3][3][16]     = A[3][3][16] ^ ((~A[4][3][16]) & A[0][3][16]);
   assign A_chi[3][3][17]     = A[3][3][17] ^ ((~A[4][3][17]) & A[0][3][17]);
   assign A_chi[3][3][18]     = A[3][3][18] ^ ((~A[4][3][18]) & A[0][3][18]);
   assign A_chi[3][3][19]     = A[3][3][19] ^ ((~A[4][3][19]) & A[0][3][19]);
   assign A_chi[3][3][20]     = A[3][3][20] ^ ((~A[4][3][20]) & A[0][3][20]);
   assign A_chi[3][3][21]     = A[3][3][21] ^ ((~A[4][3][21]) & A[0][3][21]);
   assign A_chi[3][3][22]     = A[3][3][22] ^ ((~A[4][3][22]) & A[0][3][22]);
   assign A_chi[3][3][23]     = A[3][3][23] ^ ((~A[4][3][23]) & A[0][3][23]);
   assign A_chi[3][3][24]     = A[3][3][24] ^ ((~A[4][3][24]) & A[0][3][24]);
   assign A_chi[3][3][25]     = A[3][3][25] ^ ((~A[4][3][25]) & A[0][3][25]);
   assign A_chi[3][3][26]     = A[3][3][26] ^ ((~A[4][3][26]) & A[0][3][26]);
   assign A_chi[3][3][27]     = A[3][3][27] ^ ((~A[4][3][27]) & A[0][3][27]);
   assign A_chi[3][3][28]     = A[3][3][28] ^ ((~A[4][3][28]) & A[0][3][28]);
   assign A_chi[3][3][29]     = A[3][3][29] ^ ((~A[4][3][29]) & A[0][3][29]);
   assign A_chi[3][3][30]     = A[3][3][30] ^ ((~A[4][3][30]) & A[0][3][30]);
   assign A_chi[3][3][31]     = A[3][3][31] ^ ((~A[4][3][31]) & A[0][3][31]);
   assign A_chi[3][3][32]     = A[3][3][32] ^ ((~A[4][3][32]) & A[0][3][32]);
   assign A_chi[3][3][33]     = A[3][3][33] ^ ((~A[4][3][33]) & A[0][3][33]);
   assign A_chi[3][3][34]     = A[3][3][34] ^ ((~A[4][3][34]) & A[0][3][34]);
   assign A_chi[3][3][35]     = A[3][3][35] ^ ((~A[4][3][35]) & A[0][3][35]);
   assign A_chi[3][3][36]     = A[3][3][36] ^ ((~A[4][3][36]) & A[0][3][36]);
   assign A_chi[3][3][37]     = A[3][3][37] ^ ((~A[4][3][37]) & A[0][3][37]);
   assign A_chi[3][3][38]     = A[3][3][38] ^ ((~A[4][3][38]) & A[0][3][38]);
   assign A_chi[3][3][39]     = A[3][3][39] ^ ((~A[4][3][39]) & A[0][3][39]);
   assign A_chi[3][3][40]     = A[3][3][40] ^ ((~A[4][3][40]) & A[0][3][40]);
   assign A_chi[3][3][41]     = A[3][3][41] ^ ((~A[4][3][41]) & A[0][3][41]);
   assign A_chi[3][3][42]     = A[3][3][42] ^ ((~A[4][3][42]) & A[0][3][42]);
   assign A_chi[3][3][43]     = A[3][3][43] ^ ((~A[4][3][43]) & A[0][3][43]);
   assign A_chi[3][3][44]     = A[3][3][44] ^ ((~A[4][3][44]) & A[0][3][44]);
   assign A_chi[3][3][45]     = A[3][3][45] ^ ((~A[4][3][45]) & A[0][3][45]);
   assign A_chi[3][3][46]     = A[3][3][46] ^ ((~A[4][3][46]) & A[0][3][46]);
   assign A_chi[3][3][47]     = A[3][3][47] ^ ((~A[4][3][47]) & A[0][3][47]);
   assign A_chi[3][3][48]     = A[3][3][48] ^ ((~A[4][3][48]) & A[0][3][48]);
   assign A_chi[3][3][49]     = A[3][3][49] ^ ((~A[4][3][49]) & A[0][3][49]);
   assign A_chi[3][3][50]     = A[3][3][50] ^ ((~A[4][3][50]) & A[0][3][50]);
   assign A_chi[3][3][51]     = A[3][3][51] ^ ((~A[4][3][51]) & A[0][3][51]);
   assign A_chi[3][3][52]     = A[3][3][52] ^ ((~A[4][3][52]) & A[0][3][52]);
   assign A_chi[3][3][53]     = A[3][3][53] ^ ((~A[4][3][53]) & A[0][3][53]);
   assign A_chi[3][3][54]     = A[3][3][54] ^ ((~A[4][3][54]) & A[0][3][54]);
   assign A_chi[3][3][55]     = A[3][3][55] ^ ((~A[4][3][55]) & A[0][3][55]);
   assign A_chi[3][3][56]     = A[3][3][56] ^ ((~A[4][3][56]) & A[0][3][56]);
   assign A_chi[3][3][57]     = A[3][3][57] ^ ((~A[4][3][57]) & A[0][3][57]);
   assign A_chi[3][3][58]     = A[3][3][58] ^ ((~A[4][3][58]) & A[0][3][58]);
   assign A_chi[3][3][59]     = A[3][3][59] ^ ((~A[4][3][59]) & A[0][3][59]);
   assign A_chi[3][3][60]     = A[3][3][60] ^ ((~A[4][3][60]) & A[0][3][60]);
   assign A_chi[3][3][61]     = A[3][3][61] ^ ((~A[4][3][61]) & A[0][3][61]);
   assign A_chi[3][3][62]     = A[3][3][62] ^ ((~A[4][3][62]) & A[0][3][62]);
   assign A_chi[3][3][63]     = A[3][3][63] ^ ((~A[4][3][63]) & A[0][3][63]);
   assign A_chi[3][4][0]     = A[4][3][0] ^ ((~A[0][3][0]) & A[1][3][0]);
   assign A_chi[3][4][1]     = A[4][3][1] ^ ((~A[0][3][1]) & A[1][3][1]);
   assign A_chi[3][4][2]     = A[4][3][2] ^ ((~A[0][3][2]) & A[1][3][2]);
   assign A_chi[3][4][3]     = A[4][3][3] ^ ((~A[0][3][3]) & A[1][3][3]);
   assign A_chi[3][4][4]     = A[4][3][4] ^ ((~A[0][3][4]) & A[1][3][4]);
   assign A_chi[3][4][5]     = A[4][3][5] ^ ((~A[0][3][5]) & A[1][3][5]);
   assign A_chi[3][4][6]     = A[4][3][6] ^ ((~A[0][3][6]) & A[1][3][6]);
   assign A_chi[3][4][7]     = A[4][3][7] ^ ((~A[0][3][7]) & A[1][3][7]);
   assign A_chi[3][4][8]     = A[4][3][8] ^ ((~A[0][3][8]) & A[1][3][8]);
   assign A_chi[3][4][9]     = A[4][3][9] ^ ((~A[0][3][9]) & A[1][3][9]);
   assign A_chi[3][4][10]     = A[4][3][10] ^ ((~A[0][3][10]) & A[1][3][10]);
   assign A_chi[3][4][11]     = A[4][3][11] ^ ((~A[0][3][11]) & A[1][3][11]);
   assign A_chi[3][4][12]     = A[4][3][12] ^ ((~A[0][3][12]) & A[1][3][12]);
   assign A_chi[3][4][13]     = A[4][3][13] ^ ((~A[0][3][13]) & A[1][3][13]);
   assign A_chi[3][4][14]     = A[4][3][14] ^ ((~A[0][3][14]) & A[1][3][14]);
   assign A_chi[3][4][15]     = A[4][3][15] ^ ((~A[0][3][15]) & A[1][3][15]);
   assign A_chi[3][4][16]     = A[4][3][16] ^ ((~A[0][3][16]) & A[1][3][16]);
   assign A_chi[3][4][17]     = A[4][3][17] ^ ((~A[0][3][17]) & A[1][3][17]);
   assign A_chi[3][4][18]     = A[4][3][18] ^ ((~A[0][3][18]) & A[1][3][18]);
   assign A_chi[3][4][19]     = A[4][3][19] ^ ((~A[0][3][19]) & A[1][3][19]);
   assign A_chi[3][4][20]     = A[4][3][20] ^ ((~A[0][3][20]) & A[1][3][20]);
   assign A_chi[3][4][21]     = A[4][3][21] ^ ((~A[0][3][21]) & A[1][3][21]);
   assign A_chi[3][4][22]     = A[4][3][22] ^ ((~A[0][3][22]) & A[1][3][22]);
   assign A_chi[3][4][23]     = A[4][3][23] ^ ((~A[0][3][23]) & A[1][3][23]);
   assign A_chi[3][4][24]     = A[4][3][24] ^ ((~A[0][3][24]) & A[1][3][24]);
   assign A_chi[3][4][25]     = A[4][3][25] ^ ((~A[0][3][25]) & A[1][3][25]);
   assign A_chi[3][4][26]     = A[4][3][26] ^ ((~A[0][3][26]) & A[1][3][26]);
   assign A_chi[3][4][27]     = A[4][3][27] ^ ((~A[0][3][27]) & A[1][3][27]);
   assign A_chi[3][4][28]     = A[4][3][28] ^ ((~A[0][3][28]) & A[1][3][28]);
   assign A_chi[3][4][29]     = A[4][3][29] ^ ((~A[0][3][29]) & A[1][3][29]);
   assign A_chi[3][4][30]     = A[4][3][30] ^ ((~A[0][3][30]) & A[1][3][30]);
   assign A_chi[3][4][31]     = A[4][3][31] ^ ((~A[0][3][31]) & A[1][3][31]);
   assign A_chi[3][4][32]     = A[4][3][32] ^ ((~A[0][3][32]) & A[1][3][32]);
   assign A_chi[3][4][33]     = A[4][3][33] ^ ((~A[0][3][33]) & A[1][3][33]);
   assign A_chi[3][4][34]     = A[4][3][34] ^ ((~A[0][3][34]) & A[1][3][34]);
   assign A_chi[3][4][35]     = A[4][3][35] ^ ((~A[0][3][35]) & A[1][3][35]);
   assign A_chi[3][4][36]     = A[4][3][36] ^ ((~A[0][3][36]) & A[1][3][36]);
   assign A_chi[3][4][37]     = A[4][3][37] ^ ((~A[0][3][37]) & A[1][3][37]);
   assign A_chi[3][4][38]     = A[4][3][38] ^ ((~A[0][3][38]) & A[1][3][38]);
   assign A_chi[3][4][39]     = A[4][3][39] ^ ((~A[0][3][39]) & A[1][3][39]);
   assign A_chi[3][4][40]     = A[4][3][40] ^ ((~A[0][3][40]) & A[1][3][40]);
   assign A_chi[3][4][41]     = A[4][3][41] ^ ((~A[0][3][41]) & A[1][3][41]);
   assign A_chi[3][4][42]     = A[4][3][42] ^ ((~A[0][3][42]) & A[1][3][42]);
   assign A_chi[3][4][43]     = A[4][3][43] ^ ((~A[0][3][43]) & A[1][3][43]);
   assign A_chi[3][4][44]     = A[4][3][44] ^ ((~A[0][3][44]) & A[1][3][44]);
   assign A_chi[3][4][45]     = A[4][3][45] ^ ((~A[0][3][45]) & A[1][3][45]);
   assign A_chi[3][4][46]     = A[4][3][46] ^ ((~A[0][3][46]) & A[1][3][46]);
   assign A_chi[3][4][47]     = A[4][3][47] ^ ((~A[0][3][47]) & A[1][3][47]);
   assign A_chi[3][4][48]     = A[4][3][48] ^ ((~A[0][3][48]) & A[1][3][48]);
   assign A_chi[3][4][49]     = A[4][3][49] ^ ((~A[0][3][49]) & A[1][3][49]);
   assign A_chi[3][4][50]     = A[4][3][50] ^ ((~A[0][3][50]) & A[1][3][50]);
   assign A_chi[3][4][51]     = A[4][3][51] ^ ((~A[0][3][51]) & A[1][3][51]);
   assign A_chi[3][4][52]     = A[4][3][52] ^ ((~A[0][3][52]) & A[1][3][52]);
   assign A_chi[3][4][53]     = A[4][3][53] ^ ((~A[0][3][53]) & A[1][3][53]);
   assign A_chi[3][4][54]     = A[4][3][54] ^ ((~A[0][3][54]) & A[1][3][54]);
   assign A_chi[3][4][55]     = A[4][3][55] ^ ((~A[0][3][55]) & A[1][3][55]);
   assign A_chi[3][4][56]     = A[4][3][56] ^ ((~A[0][3][56]) & A[1][3][56]);
   assign A_chi[3][4][57]     = A[4][3][57] ^ ((~A[0][3][57]) & A[1][3][57]);
   assign A_chi[3][4][58]     = A[4][3][58] ^ ((~A[0][3][58]) & A[1][3][58]);
   assign A_chi[3][4][59]     = A[4][3][59] ^ ((~A[0][3][59]) & A[1][3][59]);
   assign A_chi[3][4][60]     = A[4][3][60] ^ ((~A[0][3][60]) & A[1][3][60]);
   assign A_chi[3][4][61]     = A[4][3][61] ^ ((~A[0][3][61]) & A[1][3][61]);
   assign A_chi[3][4][62]     = A[4][3][62] ^ ((~A[0][3][62]) & A[1][3][62]);
   assign A_chi[3][4][63]     = A[4][3][63] ^ ((~A[0][3][63]) & A[1][3][63]);
   assign A_chi[4][0][0]     = A[0][4][0] ^ ((~A[1][4][0]) & A[2][4][0]);
   assign A_chi[4][0][1]     = A[0][4][1] ^ ((~A[1][4][1]) & A[2][4][1]);
   assign A_chi[4][0][2]     = A[0][4][2] ^ ((~A[1][4][2]) & A[2][4][2]);
   assign A_chi[4][0][3]     = A[0][4][3] ^ ((~A[1][4][3]) & A[2][4][3]);
   assign A_chi[4][0][4]     = A[0][4][4] ^ ((~A[1][4][4]) & A[2][4][4]);
   assign A_chi[4][0][5]     = A[0][4][5] ^ ((~A[1][4][5]) & A[2][4][5]);
   assign A_chi[4][0][6]     = A[0][4][6] ^ ((~A[1][4][6]) & A[2][4][6]);
   assign A_chi[4][0][7]     = A[0][4][7] ^ ((~A[1][4][7]) & A[2][4][7]);
   assign A_chi[4][0][8]     = A[0][4][8] ^ ((~A[1][4][8]) & A[2][4][8]);
   assign A_chi[4][0][9]     = A[0][4][9] ^ ((~A[1][4][9]) & A[2][4][9]);
   assign A_chi[4][0][10]     = A[0][4][10] ^ ((~A[1][4][10]) & A[2][4][10]);
   assign A_chi[4][0][11]     = A[0][4][11] ^ ((~A[1][4][11]) & A[2][4][11]);
   assign A_chi[4][0][12]     = A[0][4][12] ^ ((~A[1][4][12]) & A[2][4][12]);
   assign A_chi[4][0][13]     = A[0][4][13] ^ ((~A[1][4][13]) & A[2][4][13]);
   assign A_chi[4][0][14]     = A[0][4][14] ^ ((~A[1][4][14]) & A[2][4][14]);
   assign A_chi[4][0][15]     = A[0][4][15] ^ ((~A[1][4][15]) & A[2][4][15]);
   assign A_chi[4][0][16]     = A[0][4][16] ^ ((~A[1][4][16]) & A[2][4][16]);
   assign A_chi[4][0][17]     = A[0][4][17] ^ ((~A[1][4][17]) & A[2][4][17]);
   assign A_chi[4][0][18]     = A[0][4][18] ^ ((~A[1][4][18]) & A[2][4][18]);
   assign A_chi[4][0][19]     = A[0][4][19] ^ ((~A[1][4][19]) & A[2][4][19]);
   assign A_chi[4][0][20]     = A[0][4][20] ^ ((~A[1][4][20]) & A[2][4][20]);
   assign A_chi[4][0][21]     = A[0][4][21] ^ ((~A[1][4][21]) & A[2][4][21]);
   assign A_chi[4][0][22]     = A[0][4][22] ^ ((~A[1][4][22]) & A[2][4][22]);
   assign A_chi[4][0][23]     = A[0][4][23] ^ ((~A[1][4][23]) & A[2][4][23]);
   assign A_chi[4][0][24]     = A[0][4][24] ^ ((~A[1][4][24]) & A[2][4][24]);
   assign A_chi[4][0][25]     = A[0][4][25] ^ ((~A[1][4][25]) & A[2][4][25]);
   assign A_chi[4][0][26]     = A[0][4][26] ^ ((~A[1][4][26]) & A[2][4][26]);
   assign A_chi[4][0][27]     = A[0][4][27] ^ ((~A[1][4][27]) & A[2][4][27]);
   assign A_chi[4][0][28]     = A[0][4][28] ^ ((~A[1][4][28]) & A[2][4][28]);
   assign A_chi[4][0][29]     = A[0][4][29] ^ ((~A[1][4][29]) & A[2][4][29]);
   assign A_chi[4][0][30]     = A[0][4][30] ^ ((~A[1][4][30]) & A[2][4][30]);
   assign A_chi[4][0][31]     = A[0][4][31] ^ ((~A[1][4][31]) & A[2][4][31]);
   assign A_chi[4][0][32]     = A[0][4][32] ^ ((~A[1][4][32]) & A[2][4][32]);
   assign A_chi[4][0][33]     = A[0][4][33] ^ ((~A[1][4][33]) & A[2][4][33]);
   assign A_chi[4][0][34]     = A[0][4][34] ^ ((~A[1][4][34]) & A[2][4][34]);
   assign A_chi[4][0][35]     = A[0][4][35] ^ ((~A[1][4][35]) & A[2][4][35]);
   assign A_chi[4][0][36]     = A[0][4][36] ^ ((~A[1][4][36]) & A[2][4][36]);
   assign A_chi[4][0][37]     = A[0][4][37] ^ ((~A[1][4][37]) & A[2][4][37]);
   assign A_chi[4][0][38]     = A[0][4][38] ^ ((~A[1][4][38]) & A[2][4][38]);
   assign A_chi[4][0][39]     = A[0][4][39] ^ ((~A[1][4][39]) & A[2][4][39]);
   assign A_chi[4][0][40]     = A[0][4][40] ^ ((~A[1][4][40]) & A[2][4][40]);
   assign A_chi[4][0][41]     = A[0][4][41] ^ ((~A[1][4][41]) & A[2][4][41]);
   assign A_chi[4][0][42]     = A[0][4][42] ^ ((~A[1][4][42]) & A[2][4][42]);
   assign A_chi[4][0][43]     = A[0][4][43] ^ ((~A[1][4][43]) & A[2][4][43]);
   assign A_chi[4][0][44]     = A[0][4][44] ^ ((~A[1][4][44]) & A[2][4][44]);
   assign A_chi[4][0][45]     = A[0][4][45] ^ ((~A[1][4][45]) & A[2][4][45]);
   assign A_chi[4][0][46]     = A[0][4][46] ^ ((~A[1][4][46]) & A[2][4][46]);
   assign A_chi[4][0][47]     = A[0][4][47] ^ ((~A[1][4][47]) & A[2][4][47]);
   assign A_chi[4][0][48]     = A[0][4][48] ^ ((~A[1][4][48]) & A[2][4][48]);
   assign A_chi[4][0][49]     = A[0][4][49] ^ ((~A[1][4][49]) & A[2][4][49]);
   assign A_chi[4][0][50]     = A[0][4][50] ^ ((~A[1][4][50]) & A[2][4][50]);
   assign A_chi[4][0][51]     = A[0][4][51] ^ ((~A[1][4][51]) & A[2][4][51]);
   assign A_chi[4][0][52]     = A[0][4][52] ^ ((~A[1][4][52]) & A[2][4][52]);
   assign A_chi[4][0][53]     = A[0][4][53] ^ ((~A[1][4][53]) & A[2][4][53]);
   assign A_chi[4][0][54]     = A[0][4][54] ^ ((~A[1][4][54]) & A[2][4][54]);
   assign A_chi[4][0][55]     = A[0][4][55] ^ ((~A[1][4][55]) & A[2][4][55]);
   assign A_chi[4][0][56]     = A[0][4][56] ^ ((~A[1][4][56]) & A[2][4][56]);
   assign A_chi[4][0][57]     = A[0][4][57] ^ ((~A[1][4][57]) & A[2][4][57]);
   assign A_chi[4][0][58]     = A[0][4][58] ^ ((~A[1][4][58]) & A[2][4][58]);
   assign A_chi[4][0][59]     = A[0][4][59] ^ ((~A[1][4][59]) & A[2][4][59]);
   assign A_chi[4][0][60]     = A[0][4][60] ^ ((~A[1][4][60]) & A[2][4][60]);
   assign A_chi[4][0][61]     = A[0][4][61] ^ ((~A[1][4][61]) & A[2][4][61]);
   assign A_chi[4][0][62]     = A[0][4][62] ^ ((~A[1][4][62]) & A[2][4][62]);
   assign A_chi[4][0][63]     = A[0][4][63] ^ ((~A[1][4][63]) & A[2][4][63]);
   assign A_chi[4][1][0]     = A[1][4][0] ^ ((~A[2][4][0]) & A[3][4][0]);
   assign A_chi[4][1][1]     = A[1][4][1] ^ ((~A[2][4][1]) & A[3][4][1]);
   assign A_chi[4][1][2]     = A[1][4][2] ^ ((~A[2][4][2]) & A[3][4][2]);
   assign A_chi[4][1][3]     = A[1][4][3] ^ ((~A[2][4][3]) & A[3][4][3]);
   assign A_chi[4][1][4]     = A[1][4][4] ^ ((~A[2][4][4]) & A[3][4][4]);
   assign A_chi[4][1][5]     = A[1][4][5] ^ ((~A[2][4][5]) & A[3][4][5]);
   assign A_chi[4][1][6]     = A[1][4][6] ^ ((~A[2][4][6]) & A[3][4][6]);
   assign A_chi[4][1][7]     = A[1][4][7] ^ ((~A[2][4][7]) & A[3][4][7]);
   assign A_chi[4][1][8]     = A[1][4][8] ^ ((~A[2][4][8]) & A[3][4][8]);
   assign A_chi[4][1][9]     = A[1][4][9] ^ ((~A[2][4][9]) & A[3][4][9]);
   assign A_chi[4][1][10]     = A[1][4][10] ^ ((~A[2][4][10]) & A[3][4][10]);
   assign A_chi[4][1][11]     = A[1][4][11] ^ ((~A[2][4][11]) & A[3][4][11]);
   assign A_chi[4][1][12]     = A[1][4][12] ^ ((~A[2][4][12]) & A[3][4][12]);
   assign A_chi[4][1][13]     = A[1][4][13] ^ ((~A[2][4][13]) & A[3][4][13]);
   assign A_chi[4][1][14]     = A[1][4][14] ^ ((~A[2][4][14]) & A[3][4][14]);
   assign A_chi[4][1][15]     = A[1][4][15] ^ ((~A[2][4][15]) & A[3][4][15]);
   assign A_chi[4][1][16]     = A[1][4][16] ^ ((~A[2][4][16]) & A[3][4][16]);
   assign A_chi[4][1][17]     = A[1][4][17] ^ ((~A[2][4][17]) & A[3][4][17]);
   assign A_chi[4][1][18]     = A[1][4][18] ^ ((~A[2][4][18]) & A[3][4][18]);
   assign A_chi[4][1][19]     = A[1][4][19] ^ ((~A[2][4][19]) & A[3][4][19]);
   assign A_chi[4][1][20]     = A[1][4][20] ^ ((~A[2][4][20]) & A[3][4][20]);
   assign A_chi[4][1][21]     = A[1][4][21] ^ ((~A[2][4][21]) & A[3][4][21]);
   assign A_chi[4][1][22]     = A[1][4][22] ^ ((~A[2][4][22]) & A[3][4][22]);
   assign A_chi[4][1][23]     = A[1][4][23] ^ ((~A[2][4][23]) & A[3][4][23]);
   assign A_chi[4][1][24]     = A[1][4][24] ^ ((~A[2][4][24]) & A[3][4][24]);
   assign A_chi[4][1][25]     = A[1][4][25] ^ ((~A[2][4][25]) & A[3][4][25]);
   assign A_chi[4][1][26]     = A[1][4][26] ^ ((~A[2][4][26]) & A[3][4][26]);
   assign A_chi[4][1][27]     = A[1][4][27] ^ ((~A[2][4][27]) & A[3][4][27]);
   assign A_chi[4][1][28]     = A[1][4][28] ^ ((~A[2][4][28]) & A[3][4][28]);
   assign A_chi[4][1][29]     = A[1][4][29] ^ ((~A[2][4][29]) & A[3][4][29]);
   assign A_chi[4][1][30]     = A[1][4][30] ^ ((~A[2][4][30]) & A[3][4][30]);
   assign A_chi[4][1][31]     = A[1][4][31] ^ ((~A[2][4][31]) & A[3][4][31]);
   assign A_chi[4][1][32]     = A[1][4][32] ^ ((~A[2][4][32]) & A[3][4][32]);
   assign A_chi[4][1][33]     = A[1][4][33] ^ ((~A[2][4][33]) & A[3][4][33]);
   assign A_chi[4][1][34]     = A[1][4][34] ^ ((~A[2][4][34]) & A[3][4][34]);
   assign A_chi[4][1][35]     = A[1][4][35] ^ ((~A[2][4][35]) & A[3][4][35]);
   assign A_chi[4][1][36]     = A[1][4][36] ^ ((~A[2][4][36]) & A[3][4][36]);
   assign A_chi[4][1][37]     = A[1][4][37] ^ ((~A[2][4][37]) & A[3][4][37]);
   assign A_chi[4][1][38]     = A[1][4][38] ^ ((~A[2][4][38]) & A[3][4][38]);
   assign A_chi[4][1][39]     = A[1][4][39] ^ ((~A[2][4][39]) & A[3][4][39]);
   assign A_chi[4][1][40]     = A[1][4][40] ^ ((~A[2][4][40]) & A[3][4][40]);
   assign A_chi[4][1][41]     = A[1][4][41] ^ ((~A[2][4][41]) & A[3][4][41]);
   assign A_chi[4][1][42]     = A[1][4][42] ^ ((~A[2][4][42]) & A[3][4][42]);
   assign A_chi[4][1][43]     = A[1][4][43] ^ ((~A[2][4][43]) & A[3][4][43]);
   assign A_chi[4][1][44]     = A[1][4][44] ^ ((~A[2][4][44]) & A[3][4][44]);
   assign A_chi[4][1][45]     = A[1][4][45] ^ ((~A[2][4][45]) & A[3][4][45]);
   assign A_chi[4][1][46]     = A[1][4][46] ^ ((~A[2][4][46]) & A[3][4][46]);
   assign A_chi[4][1][47]     = A[1][4][47] ^ ((~A[2][4][47]) & A[3][4][47]);
   assign A_chi[4][1][48]     = A[1][4][48] ^ ((~A[2][4][48]) & A[3][4][48]);
   assign A_chi[4][1][49]     = A[1][4][49] ^ ((~A[2][4][49]) & A[3][4][49]);
   assign A_chi[4][1][50]     = A[1][4][50] ^ ((~A[2][4][50]) & A[3][4][50]);
   assign A_chi[4][1][51]     = A[1][4][51] ^ ((~A[2][4][51]) & A[3][4][51]);
   assign A_chi[4][1][52]     = A[1][4][52] ^ ((~A[2][4][52]) & A[3][4][52]);
   assign A_chi[4][1][53]     = A[1][4][53] ^ ((~A[2][4][53]) & A[3][4][53]);
   assign A_chi[4][1][54]     = A[1][4][54] ^ ((~A[2][4][54]) & A[3][4][54]);
   assign A_chi[4][1][55]     = A[1][4][55] ^ ((~A[2][4][55]) & A[3][4][55]);
   assign A_chi[4][1][56]     = A[1][4][56] ^ ((~A[2][4][56]) & A[3][4][56]);
   assign A_chi[4][1][57]     = A[1][4][57] ^ ((~A[2][4][57]) & A[3][4][57]);
   assign A_chi[4][1][58]     = A[1][4][58] ^ ((~A[2][4][58]) & A[3][4][58]);
   assign A_chi[4][1][59]     = A[1][4][59] ^ ((~A[2][4][59]) & A[3][4][59]);
   assign A_chi[4][1][60]     = A[1][4][60] ^ ((~A[2][4][60]) & A[3][4][60]);
   assign A_chi[4][1][61]     = A[1][4][61] ^ ((~A[2][4][61]) & A[3][4][61]);
   assign A_chi[4][1][62]     = A[1][4][62] ^ ((~A[2][4][62]) & A[3][4][62]);
   assign A_chi[4][1][63]     = A[1][4][63] ^ ((~A[2][4][63]) & A[3][4][63]);
   assign A_chi[4][2][0]     = A[2][4][0] ^ ((~A[3][4][0]) & A[4][4][0]);
   assign A_chi[4][2][1]     = A[2][4][1] ^ ((~A[3][4][1]) & A[4][4][1]);
   assign A_chi[4][2][2]     = A[2][4][2] ^ ((~A[3][4][2]) & A[4][4][2]);
   assign A_chi[4][2][3]     = A[2][4][3] ^ ((~A[3][4][3]) & A[4][4][3]);
   assign A_chi[4][2][4]     = A[2][4][4] ^ ((~A[3][4][4]) & A[4][4][4]);
   assign A_chi[4][2][5]     = A[2][4][5] ^ ((~A[3][4][5]) & A[4][4][5]);
   assign A_chi[4][2][6]     = A[2][4][6] ^ ((~A[3][4][6]) & A[4][4][6]);
   assign A_chi[4][2][7]     = A[2][4][7] ^ ((~A[3][4][7]) & A[4][4][7]);
   assign A_chi[4][2][8]     = A[2][4][8] ^ ((~A[3][4][8]) & A[4][4][8]);
   assign A_chi[4][2][9]     = A[2][4][9] ^ ((~A[3][4][9]) & A[4][4][9]);
   assign A_chi[4][2][10]     = A[2][4][10] ^ ((~A[3][4][10]) & A[4][4][10]);
   assign A_chi[4][2][11]     = A[2][4][11] ^ ((~A[3][4][11]) & A[4][4][11]);
   assign A_chi[4][2][12]     = A[2][4][12] ^ ((~A[3][4][12]) & A[4][4][12]);
   assign A_chi[4][2][13]     = A[2][4][13] ^ ((~A[3][4][13]) & A[4][4][13]);
   assign A_chi[4][2][14]     = A[2][4][14] ^ ((~A[3][4][14]) & A[4][4][14]);
   assign A_chi[4][2][15]     = A[2][4][15] ^ ((~A[3][4][15]) & A[4][4][15]);
   assign A_chi[4][2][16]     = A[2][4][16] ^ ((~A[3][4][16]) & A[4][4][16]);
   assign A_chi[4][2][17]     = A[2][4][17] ^ ((~A[3][4][17]) & A[4][4][17]);
   assign A_chi[4][2][18]     = A[2][4][18] ^ ((~A[3][4][18]) & A[4][4][18]);
   assign A_chi[4][2][19]     = A[2][4][19] ^ ((~A[3][4][19]) & A[4][4][19]);
   assign A_chi[4][2][20]     = A[2][4][20] ^ ((~A[3][4][20]) & A[4][4][20]);
   assign A_chi[4][2][21]     = A[2][4][21] ^ ((~A[3][4][21]) & A[4][4][21]);
   assign A_chi[4][2][22]     = A[2][4][22] ^ ((~A[3][4][22]) & A[4][4][22]);
   assign A_chi[4][2][23]     = A[2][4][23] ^ ((~A[3][4][23]) & A[4][4][23]);
   assign A_chi[4][2][24]     = A[2][4][24] ^ ((~A[3][4][24]) & A[4][4][24]);
   assign A_chi[4][2][25]     = A[2][4][25] ^ ((~A[3][4][25]) & A[4][4][25]);
   assign A_chi[4][2][26]     = A[2][4][26] ^ ((~A[3][4][26]) & A[4][4][26]);
   assign A_chi[4][2][27]     = A[2][4][27] ^ ((~A[3][4][27]) & A[4][4][27]);
   assign A_chi[4][2][28]     = A[2][4][28] ^ ((~A[3][4][28]) & A[4][4][28]);
   assign A_chi[4][2][29]     = A[2][4][29] ^ ((~A[3][4][29]) & A[4][4][29]);
   assign A_chi[4][2][30]     = A[2][4][30] ^ ((~A[3][4][30]) & A[4][4][30]);
   assign A_chi[4][2][31]     = A[2][4][31] ^ ((~A[3][4][31]) & A[4][4][31]);
   assign A_chi[4][2][32]     = A[2][4][32] ^ ((~A[3][4][32]) & A[4][4][32]);
   assign A_chi[4][2][33]     = A[2][4][33] ^ ((~A[3][4][33]) & A[4][4][33]);
   assign A_chi[4][2][34]     = A[2][4][34] ^ ((~A[3][4][34]) & A[4][4][34]);
   assign A_chi[4][2][35]     = A[2][4][35] ^ ((~A[3][4][35]) & A[4][4][35]);
   assign A_chi[4][2][36]     = A[2][4][36] ^ ((~A[3][4][36]) & A[4][4][36]);
   assign A_chi[4][2][37]     = A[2][4][37] ^ ((~A[3][4][37]) & A[4][4][37]);
   assign A_chi[4][2][38]     = A[2][4][38] ^ ((~A[3][4][38]) & A[4][4][38]);
   assign A_chi[4][2][39]     = A[2][4][39] ^ ((~A[3][4][39]) & A[4][4][39]);
   assign A_chi[4][2][40]     = A[2][4][40] ^ ((~A[3][4][40]) & A[4][4][40]);
   assign A_chi[4][2][41]     = A[2][4][41] ^ ((~A[3][4][41]) & A[4][4][41]);
   assign A_chi[4][2][42]     = A[2][4][42] ^ ((~A[3][4][42]) & A[4][4][42]);
   assign A_chi[4][2][43]     = A[2][4][43] ^ ((~A[3][4][43]) & A[4][4][43]);
   assign A_chi[4][2][44]     = A[2][4][44] ^ ((~A[3][4][44]) & A[4][4][44]);
   assign A_chi[4][2][45]     = A[2][4][45] ^ ((~A[3][4][45]) & A[4][4][45]);
   assign A_chi[4][2][46]     = A[2][4][46] ^ ((~A[3][4][46]) & A[4][4][46]);
   assign A_chi[4][2][47]     = A[2][4][47] ^ ((~A[3][4][47]) & A[4][4][47]);
   assign A_chi[4][2][48]     = A[2][4][48] ^ ((~A[3][4][48]) & A[4][4][48]);
   assign A_chi[4][2][49]     = A[2][4][49] ^ ((~A[3][4][49]) & A[4][4][49]);
   assign A_chi[4][2][50]     = A[2][4][50] ^ ((~A[3][4][50]) & A[4][4][50]);
   assign A_chi[4][2][51]     = A[2][4][51] ^ ((~A[3][4][51]) & A[4][4][51]);
   assign A_chi[4][2][52]     = A[2][4][52] ^ ((~A[3][4][52]) & A[4][4][52]);
   assign A_chi[4][2][53]     = A[2][4][53] ^ ((~A[3][4][53]) & A[4][4][53]);
   assign A_chi[4][2][54]     = A[2][4][54] ^ ((~A[3][4][54]) & A[4][4][54]);
   assign A_chi[4][2][55]     = A[2][4][55] ^ ((~A[3][4][55]) & A[4][4][55]);
   assign A_chi[4][2][56]     = A[2][4][56] ^ ((~A[3][4][56]) & A[4][4][56]);
   assign A_chi[4][2][57]     = A[2][4][57] ^ ((~A[3][4][57]) & A[4][4][57]);
   assign A_chi[4][2][58]     = A[2][4][58] ^ ((~A[3][4][58]) & A[4][4][58]);
   assign A_chi[4][2][59]     = A[2][4][59] ^ ((~A[3][4][59]) & A[4][4][59]);
   assign A_chi[4][2][60]     = A[2][4][60] ^ ((~A[3][4][60]) & A[4][4][60]);
   assign A_chi[4][2][61]     = A[2][4][61] ^ ((~A[3][4][61]) & A[4][4][61]);
   assign A_chi[4][2][62]     = A[2][4][62] ^ ((~A[3][4][62]) & A[4][4][62]);
   assign A_chi[4][2][63]     = A[2][4][63] ^ ((~A[3][4][63]) & A[4][4][63]);
   assign A_chi[4][3][0]     = A[3][4][0] ^ ((~A[4][4][0]) & A[0][4][0]);
   assign A_chi[4][3][1]     = A[3][4][1] ^ ((~A[4][4][1]) & A[0][4][1]);
   assign A_chi[4][3][2]     = A[3][4][2] ^ ((~A[4][4][2]) & A[0][4][2]);
   assign A_chi[4][3][3]     = A[3][4][3] ^ ((~A[4][4][3]) & A[0][4][3]);
   assign A_chi[4][3][4]     = A[3][4][4] ^ ((~A[4][4][4]) & A[0][4][4]);
   assign A_chi[4][3][5]     = A[3][4][5] ^ ((~A[4][4][5]) & A[0][4][5]);
   assign A_chi[4][3][6]     = A[3][4][6] ^ ((~A[4][4][6]) & A[0][4][6]);
   assign A_chi[4][3][7]     = A[3][4][7] ^ ((~A[4][4][7]) & A[0][4][7]);
   assign A_chi[4][3][8]     = A[3][4][8] ^ ((~A[4][4][8]) & A[0][4][8]);
   assign A_chi[4][3][9]     = A[3][4][9] ^ ((~A[4][4][9]) & A[0][4][9]);
   assign A_chi[4][3][10]     = A[3][4][10] ^ ((~A[4][4][10]) & A[0][4][10]);
   assign A_chi[4][3][11]     = A[3][4][11] ^ ((~A[4][4][11]) & A[0][4][11]);
   assign A_chi[4][3][12]     = A[3][4][12] ^ ((~A[4][4][12]) & A[0][4][12]);
   assign A_chi[4][3][13]     = A[3][4][13] ^ ((~A[4][4][13]) & A[0][4][13]);
   assign A_chi[4][3][14]     = A[3][4][14] ^ ((~A[4][4][14]) & A[0][4][14]);
   assign A_chi[4][3][15]     = A[3][4][15] ^ ((~A[4][4][15]) & A[0][4][15]);
   assign A_chi[4][3][16]     = A[3][4][16] ^ ((~A[4][4][16]) & A[0][4][16]);
   assign A_chi[4][3][17]     = A[3][4][17] ^ ((~A[4][4][17]) & A[0][4][17]);
   assign A_chi[4][3][18]     = A[3][4][18] ^ ((~A[4][4][18]) & A[0][4][18]);
   assign A_chi[4][3][19]     = A[3][4][19] ^ ((~A[4][4][19]) & A[0][4][19]);
   assign A_chi[4][3][20]     = A[3][4][20] ^ ((~A[4][4][20]) & A[0][4][20]);
   assign A_chi[4][3][21]     = A[3][4][21] ^ ((~A[4][4][21]) & A[0][4][21]);
   assign A_chi[4][3][22]     = A[3][4][22] ^ ((~A[4][4][22]) & A[0][4][22]);
   assign A_chi[4][3][23]     = A[3][4][23] ^ ((~A[4][4][23]) & A[0][4][23]);
   assign A_chi[4][3][24]     = A[3][4][24] ^ ((~A[4][4][24]) & A[0][4][24]);
   assign A_chi[4][3][25]     = A[3][4][25] ^ ((~A[4][4][25]) & A[0][4][25]);
   assign A_chi[4][3][26]     = A[3][4][26] ^ ((~A[4][4][26]) & A[0][4][26]);
   assign A_chi[4][3][27]     = A[3][4][27] ^ ((~A[4][4][27]) & A[0][4][27]);
   assign A_chi[4][3][28]     = A[3][4][28] ^ ((~A[4][4][28]) & A[0][4][28]);
   assign A_chi[4][3][29]     = A[3][4][29] ^ ((~A[4][4][29]) & A[0][4][29]);
   assign A_chi[4][3][30]     = A[3][4][30] ^ ((~A[4][4][30]) & A[0][4][30]);
   assign A_chi[4][3][31]     = A[3][4][31] ^ ((~A[4][4][31]) & A[0][4][31]);
   assign A_chi[4][3][32]     = A[3][4][32] ^ ((~A[4][4][32]) & A[0][4][32]);
   assign A_chi[4][3][33]     = A[3][4][33] ^ ((~A[4][4][33]) & A[0][4][33]);
   assign A_chi[4][3][34]     = A[3][4][34] ^ ((~A[4][4][34]) & A[0][4][34]);
   assign A_chi[4][3][35]     = A[3][4][35] ^ ((~A[4][4][35]) & A[0][4][35]);
   assign A_chi[4][3][36]     = A[3][4][36] ^ ((~A[4][4][36]) & A[0][4][36]);
   assign A_chi[4][3][37]     = A[3][4][37] ^ ((~A[4][4][37]) & A[0][4][37]);
   assign A_chi[4][3][38]     = A[3][4][38] ^ ((~A[4][4][38]) & A[0][4][38]);
   assign A_chi[4][3][39]     = A[3][4][39] ^ ((~A[4][4][39]) & A[0][4][39]);
   assign A_chi[4][3][40]     = A[3][4][40] ^ ((~A[4][4][40]) & A[0][4][40]);
   assign A_chi[4][3][41]     = A[3][4][41] ^ ((~A[4][4][41]) & A[0][4][41]);
   assign A_chi[4][3][42]     = A[3][4][42] ^ ((~A[4][4][42]) & A[0][4][42]);
   assign A_chi[4][3][43]     = A[3][4][43] ^ ((~A[4][4][43]) & A[0][4][43]);
   assign A_chi[4][3][44]     = A[3][4][44] ^ ((~A[4][4][44]) & A[0][4][44]);
   assign A_chi[4][3][45]     = A[3][4][45] ^ ((~A[4][4][45]) & A[0][4][45]);
   assign A_chi[4][3][46]     = A[3][4][46] ^ ((~A[4][4][46]) & A[0][4][46]);
   assign A_chi[4][3][47]     = A[3][4][47] ^ ((~A[4][4][47]) & A[0][4][47]);
   assign A_chi[4][3][48]     = A[3][4][48] ^ ((~A[4][4][48]) & A[0][4][48]);
   assign A_chi[4][3][49]     = A[3][4][49] ^ ((~A[4][4][49]) & A[0][4][49]);
   assign A_chi[4][3][50]     = A[3][4][50] ^ ((~A[4][4][50]) & A[0][4][50]);
   assign A_chi[4][3][51]     = A[3][4][51] ^ ((~A[4][4][51]) & A[0][4][51]);
   assign A_chi[4][3][52]     = A[3][4][52] ^ ((~A[4][4][52]) & A[0][4][52]);
   assign A_chi[4][3][53]     = A[3][4][53] ^ ((~A[4][4][53]) & A[0][4][53]);
   assign A_chi[4][3][54]     = A[3][4][54] ^ ((~A[4][4][54]) & A[0][4][54]);
   assign A_chi[4][3][55]     = A[3][4][55] ^ ((~A[4][4][55]) & A[0][4][55]);
   assign A_chi[4][3][56]     = A[3][4][56] ^ ((~A[4][4][56]) & A[0][4][56]);
   assign A_chi[4][3][57]     = A[3][4][57] ^ ((~A[4][4][57]) & A[0][4][57]);
   assign A_chi[4][3][58]     = A[3][4][58] ^ ((~A[4][4][58]) & A[0][4][58]);
   assign A_chi[4][3][59]     = A[3][4][59] ^ ((~A[4][4][59]) & A[0][4][59]);
   assign A_chi[4][3][60]     = A[3][4][60] ^ ((~A[4][4][60]) & A[0][4][60]);
   assign A_chi[4][3][61]     = A[3][4][61] ^ ((~A[4][4][61]) & A[0][4][61]);
   assign A_chi[4][3][62]     = A[3][4][62] ^ ((~A[4][4][62]) & A[0][4][62]);
   assign A_chi[4][3][63]     = A[3][4][63] ^ ((~A[4][4][63]) & A[0][4][63]);
   assign A_chi[4][4][0]     = A[4][4][0] ^ ((~A[0][4][0]) & A[1][4][0]);
   assign A_chi[4][4][1]     = A[4][4][1] ^ ((~A[0][4][1]) & A[1][4][1]);
   assign A_chi[4][4][2]     = A[4][4][2] ^ ((~A[0][4][2]) & A[1][4][2]);
   assign A_chi[4][4][3]     = A[4][4][3] ^ ((~A[0][4][3]) & A[1][4][3]);
   assign A_chi[4][4][4]     = A[4][4][4] ^ ((~A[0][4][4]) & A[1][4][4]);
   assign A_chi[4][4][5]     = A[4][4][5] ^ ((~A[0][4][5]) & A[1][4][5]);
   assign A_chi[4][4][6]     = A[4][4][6] ^ ((~A[0][4][6]) & A[1][4][6]);
   assign A_chi[4][4][7]     = A[4][4][7] ^ ((~A[0][4][7]) & A[1][4][7]);
   assign A_chi[4][4][8]     = A[4][4][8] ^ ((~A[0][4][8]) & A[1][4][8]);
   assign A_chi[4][4][9]     = A[4][4][9] ^ ((~A[0][4][9]) & A[1][4][9]);
   assign A_chi[4][4][10]     = A[4][4][10] ^ ((~A[0][4][10]) & A[1][4][10]);
   assign A_chi[4][4][11]     = A[4][4][11] ^ ((~A[0][4][11]) & A[1][4][11]);
   assign A_chi[4][4][12]     = A[4][4][12] ^ ((~A[0][4][12]) & A[1][4][12]);
   assign A_chi[4][4][13]     = A[4][4][13] ^ ((~A[0][4][13]) & A[1][4][13]);
   assign A_chi[4][4][14]     = A[4][4][14] ^ ((~A[0][4][14]) & A[1][4][14]);
   assign A_chi[4][4][15]     = A[4][4][15] ^ ((~A[0][4][15]) & A[1][4][15]);
   assign A_chi[4][4][16]     = A[4][4][16] ^ ((~A[0][4][16]) & A[1][4][16]);
   assign A_chi[4][4][17]     = A[4][4][17] ^ ((~A[0][4][17]) & A[1][4][17]);
   assign A_chi[4][4][18]     = A[4][4][18] ^ ((~A[0][4][18]) & A[1][4][18]);
   assign A_chi[4][4][19]     = A[4][4][19] ^ ((~A[0][4][19]) & A[1][4][19]);
   assign A_chi[4][4][20]     = A[4][4][20] ^ ((~A[0][4][20]) & A[1][4][20]);
   assign A_chi[4][4][21]     = A[4][4][21] ^ ((~A[0][4][21]) & A[1][4][21]);
   assign A_chi[4][4][22]     = A[4][4][22] ^ ((~A[0][4][22]) & A[1][4][22]);
   assign A_chi[4][4][23]     = A[4][4][23] ^ ((~A[0][4][23]) & A[1][4][23]);
   assign A_chi[4][4][24]     = A[4][4][24] ^ ((~A[0][4][24]) & A[1][4][24]);
   assign A_chi[4][4][25]     = A[4][4][25] ^ ((~A[0][4][25]) & A[1][4][25]);
   assign A_chi[4][4][26]     = A[4][4][26] ^ ((~A[0][4][26]) & A[1][4][26]);
   assign A_chi[4][4][27]     = A[4][4][27] ^ ((~A[0][4][27]) & A[1][4][27]);
   assign A_chi[4][4][28]     = A[4][4][28] ^ ((~A[0][4][28]) & A[1][4][28]);
   assign A_chi[4][4][29]     = A[4][4][29] ^ ((~A[0][4][29]) & A[1][4][29]);
   assign A_chi[4][4][30]     = A[4][4][30] ^ ((~A[0][4][30]) & A[1][4][30]);
   assign A_chi[4][4][31]     = A[4][4][31] ^ ((~A[0][4][31]) & A[1][4][31]);
   assign A_chi[4][4][32]     = A[4][4][32] ^ ((~A[0][4][32]) & A[1][4][32]);
   assign A_chi[4][4][33]     = A[4][4][33] ^ ((~A[0][4][33]) & A[1][4][33]);
   assign A_chi[4][4][34]     = A[4][4][34] ^ ((~A[0][4][34]) & A[1][4][34]);
   assign A_chi[4][4][35]     = A[4][4][35] ^ ((~A[0][4][35]) & A[1][4][35]);
   assign A_chi[4][4][36]     = A[4][4][36] ^ ((~A[0][4][36]) & A[1][4][36]);
   assign A_chi[4][4][37]     = A[4][4][37] ^ ((~A[0][4][37]) & A[1][4][37]);
   assign A_chi[4][4][38]     = A[4][4][38] ^ ((~A[0][4][38]) & A[1][4][38]);
   assign A_chi[4][4][39]     = A[4][4][39] ^ ((~A[0][4][39]) & A[1][4][39]);
   assign A_chi[4][4][40]     = A[4][4][40] ^ ((~A[0][4][40]) & A[1][4][40]);
   assign A_chi[4][4][41]     = A[4][4][41] ^ ((~A[0][4][41]) & A[1][4][41]);
   assign A_chi[4][4][42]     = A[4][4][42] ^ ((~A[0][4][42]) & A[1][4][42]);
   assign A_chi[4][4][43]     = A[4][4][43] ^ ((~A[0][4][43]) & A[1][4][43]);
   assign A_chi[4][4][44]     = A[4][4][44] ^ ((~A[0][4][44]) & A[1][4][44]);
   assign A_chi[4][4][45]     = A[4][4][45] ^ ((~A[0][4][45]) & A[1][4][45]);
   assign A_chi[4][4][46]     = A[4][4][46] ^ ((~A[0][4][46]) & A[1][4][46]);
   assign A_chi[4][4][47]     = A[4][4][47] ^ ((~A[0][4][47]) & A[1][4][47]);
   assign A_chi[4][4][48]     = A[4][4][48] ^ ((~A[0][4][48]) & A[1][4][48]);
   assign A_chi[4][4][49]     = A[4][4][49] ^ ((~A[0][4][49]) & A[1][4][49]);
   assign A_chi[4][4][50]     = A[4][4][50] ^ ((~A[0][4][50]) & A[1][4][50]);
   assign A_chi[4][4][51]     = A[4][4][51] ^ ((~A[0][4][51]) & A[1][4][51]);
   assign A_chi[4][4][52]     = A[4][4][52] ^ ((~A[0][4][52]) & A[1][4][52]);
   assign A_chi[4][4][53]     = A[4][4][53] ^ ((~A[0][4][53]) & A[1][4][53]);
   assign A_chi[4][4][54]     = A[4][4][54] ^ ((~A[0][4][54]) & A[1][4][54]);
   assign A_chi[4][4][55]     = A[4][4][55] ^ ((~A[0][4][55]) & A[1][4][55]);
   assign A_chi[4][4][56]     = A[4][4][56] ^ ((~A[0][4][56]) & A[1][4][56]);
   assign A_chi[4][4][57]     = A[4][4][57] ^ ((~A[0][4][57]) & A[1][4][57]);
   assign A_chi[4][4][58]     = A[4][4][58] ^ ((~A[0][4][58]) & A[1][4][58]);
   assign A_chi[4][4][59]     = A[4][4][59] ^ ((~A[0][4][59]) & A[1][4][59]);
   assign A_chi[4][4][60]     = A[4][4][60] ^ ((~A[0][4][60]) & A[1][4][60]);
   assign A_chi[4][4][61]     = A[4][4][61] ^ ((~A[0][4][61]) & A[1][4][61]);
   assign A_chi[4][4][62]     = A[4][4][62] ^ ((~A[0][4][62]) & A[1][4][62]);
   assign A_chi[4][4][63]     = A[4][4][63] ^ ((~A[0][4][63]) & A[1][4][63]);
//--------------------------- IOTA ---------------------------

    // Define round constants
    reg [63:0] RC;
    always @(*) begin
        case (round_index)
            5'd0: RC   = 64'h0000000000000001;
            5'd1: RC   = 64'h0000000000008082;
            5'd2: RC   = 64'h800000000000808A;
            5'd3: RC   = 64'h8000000080008000;
            5'd4: RC   = 64'h000000000000808B;
            5'd5: RC   = 64'h0000000080000001;
            5'd6: RC   = 64'h8000000080008081;
            5'd7: RC   = 64'h8000000000008009;
            5'd8: RC   = 64'h000000000000008A;
            5'd9: RC   = 64'h0000000000000088;
            5'd10: RC   = 64'h0000000080008009;
            5'd11: RC   = 64'h000000008000000A;
            5'd12: RC   = 64'h000000008000808B;
            5'd13: RC   = 64'h800000000000008B;
            5'd14: RC   = 64'h8000000000008089;
            5'd15: RC   = 64'h8000000000008003;
            5'd16: RC   = 64'h8000000000008002;
            5'd17: RC   = 64'h8000000000000080;
            5'd18: RC   = 64'h000000000000800A;
            5'd19: RC   = 64'h800000008000000A;
            5'd20: RC   = 64'h8000000080008081;
            5'd21: RC   = 64'h8000000000008080;
            5'd22: RC   = 64'h0000000080000001;
            5'd23: RC   = 64'h8000000080008008;
            default: RC = 64'h0;
        endcase
    end

    // Apply Iota step
    always @(*) begin
        A_iota[0][0] = A[0][0];
        A_iota[1][0] = A[1][0];
        A_iota[2][0] = A[2][0];
        A_iota[3][0] = A[3][0];
        A_iota[4][0] = A[4][0];
        A_iota[0][1] = A[0][1];
        A_iota[1][1] = A[1][1];
        A_iota[2][1] = A[2][1];
        A_iota[3][1] = A[3][1];
        A_iota[4][1] = A[4][1];
        A_iota[0][2] = A[0][2];
        A_iota[1][2] = A[1][2];
        A_iota[2][2] = A[2][2];
        A_iota[3][2] = A[3][2];
        A_iota[4][2] = A[4][2];
        A_iota[0][3] = A[0][3];
        A_iota[1][3] = A[1][3];
        A_iota[2][3] = A[2][3];
        A_iota[3][3] = A[3][3];
        A_iota[4][3] = A[4][3];
        A_iota[0][4] = A[0][4];
        A_iota[1][4] = A[1][4];
        A_iota[2][4] = A[2][4];
        A_iota[3][4] = A[3][4];
        A_iota[4][4] = A[4][4];
        A_iota[0][0]  = A[0][0] ^ RC;  // XOR RC with A[0][0]
    end

    // Deflatten 3D array into S_out
    assign S_out[0]  = A_iota[0][0][0];
    assign S_out[64]  = A_iota[1][0][0];
    assign S_out[128]  = A_iota[2][0][0];
    assign S_out[192]  = A_iota[3][0][0];
    assign S_out[256]  = A_iota[4][0][0];
    assign S_out[320]  = A_iota[0][1][0];
    assign S_out[384]  = A_iota[1][1][0];
    assign S_out[448]  = A_iota[2][1][0];
    assign S_out[512]  = A_iota[3][1][0];
    assign S_out[576]  = A_iota[4][1][0];
    assign S_out[640]  = A_iota[0][2][0];
    assign S_out[704]  = A_iota[1][2][0];
    assign S_out[768]  = A_iota[2][2][0];
    assign S_out[832]  = A_iota[3][2][0];
    assign S_out[896]  = A_iota[4][2][0];
    assign S_out[960]  = A_iota[0][3][0];
    assign S_out[1024]  = A_iota[1][3][0];
    assign S_out[1088]  = A_iota[2][3][0];
    assign S_out[1152]  = A_iota[3][3][0];
    assign S_out[1216]  = A_iota[4][3][0];
    assign S_out[1280]  = A_iota[0][4][0];
    assign S_out[1344]  = A_iota[1][4][0];
    assign S_out[1408]  = A_iota[2][4][0];
    assign S_out[1472]  = A_iota[3][4][0];
    assign S_out[1536]  = A_iota[4][4][0];
    assign S_out[1]  = A_iota[0][0][1];
    assign S_out[65]  = A_iota[1][0][1];
    assign S_out[129]  = A_iota[2][0][1];
    assign S_out[193]  = A_iota[3][0][1];
    assign S_out[257]  = A_iota[4][0][1];
    assign S_out[321]  = A_iota[0][1][1];
    assign S_out[385]  = A_iota[1][1][1];
    assign S_out[449]  = A_iota[2][1][1];
    assign S_out[513]  = A_iota[3][1][1];
    assign S_out[577]  = A_iota[4][1][1];
    assign S_out[641]  = A_iota[0][2][1];
    assign S_out[705]  = A_iota[1][2][1];
    assign S_out[769]  = A_iota[2][2][1];
    assign S_out[833]  = A_iota[3][2][1];
    assign S_out[897]  = A_iota[4][2][1];
    assign S_out[961]  = A_iota[0][3][1];
    assign S_out[1025]  = A_iota[1][3][1];
    assign S_out[1089]  = A_iota[2][3][1];
    assign S_out[1153]  = A_iota[3][3][1];
    assign S_out[1217]  = A_iota[4][3][1];
    assign S_out[1281]  = A_iota[0][4][1];
    assign S_out[1345]  = A_iota[1][4][1];
    assign S_out[1409]  = A_iota[2][4][1];
    assign S_out[1473]  = A_iota[3][4][1];
    assign S_out[1537]  = A_iota[4][4][1];
    assign S_out[2]  = A_iota[0][0][2];
    assign S_out[66]  = A_iota[1][0][2];
    assign S_out[130]  = A_iota[2][0][2];
    assign S_out[194]  = A_iota[3][0][2];
    assign S_out[258]  = A_iota[4][0][2];
    assign S_out[322]  = A_iota[0][1][2];
    assign S_out[386]  = A_iota[1][1][2];
    assign S_out[450]  = A_iota[2][1][2];
    assign S_out[514]  = A_iota[3][1][2];
    assign S_out[578]  = A_iota[4][1][2];
    assign S_out[642]  = A_iota[0][2][2];
    assign S_out[706]  = A_iota[1][2][2];
    assign S_out[770]  = A_iota[2][2][2];
    assign S_out[834]  = A_iota[3][2][2];
    assign S_out[898]  = A_iota[4][2][2];
    assign S_out[962]  = A_iota[0][3][2];
    assign S_out[1026]  = A_iota[1][3][2];
    assign S_out[1090]  = A_iota[2][3][2];
    assign S_out[1154]  = A_iota[3][3][2];
    assign S_out[1218]  = A_iota[4][3][2];
    assign S_out[1282]  = A_iota[0][4][2];
    assign S_out[1346]  = A_iota[1][4][2];
    assign S_out[1410]  = A_iota[2][4][2];
    assign S_out[1474]  = A_iota[3][4][2];
    assign S_out[1538]  = A_iota[4][4][2];
    assign S_out[3]  = A_iota[0][0][3];
    assign S_out[67]  = A_iota[1][0][3];
    assign S_out[131]  = A_iota[2][0][3];
    assign S_out[195]  = A_iota[3][0][3];
    assign S_out[259]  = A_iota[4][0][3];
    assign S_out[323]  = A_iota[0][1][3];
    assign S_out[387]  = A_iota[1][1][3];
    assign S_out[451]  = A_iota[2][1][3];
    assign S_out[515]  = A_iota[3][1][3];
    assign S_out[579]  = A_iota[4][1][3];
    assign S_out[643]  = A_iota[0][2][3];
    assign S_out[707]  = A_iota[1][2][3];
    assign S_out[771]  = A_iota[2][2][3];
    assign S_out[835]  = A_iota[3][2][3];
    assign S_out[899]  = A_iota[4][2][3];
    assign S_out[963]  = A_iota[0][3][3];
    assign S_out[1027]  = A_iota[1][3][3];
    assign S_out[1091]  = A_iota[2][3][3];
    assign S_out[1155]  = A_iota[3][3][3];
    assign S_out[1219]  = A_iota[4][3][3];
    assign S_out[1283]  = A_iota[0][4][3];
    assign S_out[1347]  = A_iota[1][4][3];
    assign S_out[1411]  = A_iota[2][4][3];
    assign S_out[1475]  = A_iota[3][4][3];
    assign S_out[1539]  = A_iota[4][4][3];
    assign S_out[4]  = A_iota[0][0][4];
    assign S_out[68]  = A_iota[1][0][4];
    assign S_out[132]  = A_iota[2][0][4];
    assign S_out[196]  = A_iota[3][0][4];
    assign S_out[260]  = A_iota[4][0][4];
    assign S_out[324]  = A_iota[0][1][4];
    assign S_out[388]  = A_iota[1][1][4];
    assign S_out[452]  = A_iota[2][1][4];
    assign S_out[516]  = A_iota[3][1][4];
    assign S_out[580]  = A_iota[4][1][4];
    assign S_out[644]  = A_iota[0][2][4];
    assign S_out[708]  = A_iota[1][2][4];
    assign S_out[772]  = A_iota[2][2][4];
    assign S_out[836]  = A_iota[3][2][4];
    assign S_out[900]  = A_iota[4][2][4];
    assign S_out[964]  = A_iota[0][3][4];
    assign S_out[1028]  = A_iota[1][3][4];
    assign S_out[1092]  = A_iota[2][3][4];
    assign S_out[1156]  = A_iota[3][3][4];
    assign S_out[1220]  = A_iota[4][3][4];
    assign S_out[1284]  = A_iota[0][4][4];
    assign S_out[1348]  = A_iota[1][4][4];
    assign S_out[1412]  = A_iota[2][4][4];
    assign S_out[1476]  = A_iota[3][4][4];
    assign S_out[1540]  = A_iota[4][4][4];
    assign S_out[5]  = A_iota[0][0][5];
    assign S_out[69]  = A_iota[1][0][5];
    assign S_out[133]  = A_iota[2][0][5];
    assign S_out[197]  = A_iota[3][0][5];
    assign S_out[261]  = A_iota[4][0][5];
    assign S_out[325]  = A_iota[0][1][5];
    assign S_out[389]  = A_iota[1][1][5];
    assign S_out[453]  = A_iota[2][1][5];
    assign S_out[517]  = A_iota[3][1][5];
    assign S_out[581]  = A_iota[4][1][5];
    assign S_out[645]  = A_iota[0][2][5];
    assign S_out[709]  = A_iota[1][2][5];
    assign S_out[773]  = A_iota[2][2][5];
    assign S_out[837]  = A_iota[3][2][5];
    assign S_out[901]  = A_iota[4][2][5];
    assign S_out[965]  = A_iota[0][3][5];
    assign S_out[1029]  = A_iota[1][3][5];
    assign S_out[1093]  = A_iota[2][3][5];
    assign S_out[1157]  = A_iota[3][3][5];
    assign S_out[1221]  = A_iota[4][3][5];
    assign S_out[1285]  = A_iota[0][4][5];
    assign S_out[1349]  = A_iota[1][4][5];
    assign S_out[1413]  = A_iota[2][4][5];
    assign S_out[1477]  = A_iota[3][4][5];
    assign S_out[1541]  = A_iota[4][4][5];
    assign S_out[6]  = A_iota[0][0][6];
    assign S_out[70]  = A_iota[1][0][6];
    assign S_out[134]  = A_iota[2][0][6];
    assign S_out[198]  = A_iota[3][0][6];
    assign S_out[262]  = A_iota[4][0][6];
    assign S_out[326]  = A_iota[0][1][6];
    assign S_out[390]  = A_iota[1][1][6];
    assign S_out[454]  = A_iota[2][1][6];
    assign S_out[518]  = A_iota[3][1][6];
    assign S_out[582]  = A_iota[4][1][6];
    assign S_out[646]  = A_iota[0][2][6];
    assign S_out[710]  = A_iota[1][2][6];
    assign S_out[774]  = A_iota[2][2][6];
    assign S_out[838]  = A_iota[3][2][6];
    assign S_out[902]  = A_iota[4][2][6];
    assign S_out[966]  = A_iota[0][3][6];
    assign S_out[1030]  = A_iota[1][3][6];
    assign S_out[1094]  = A_iota[2][3][6];
    assign S_out[1158]  = A_iota[3][3][6];
    assign S_out[1222]  = A_iota[4][3][6];
    assign S_out[1286]  = A_iota[0][4][6];
    assign S_out[1350]  = A_iota[1][4][6];
    assign S_out[1414]  = A_iota[2][4][6];
    assign S_out[1478]  = A_iota[3][4][6];
    assign S_out[1542]  = A_iota[4][4][6];
    assign S_out[7]  = A_iota[0][0][7];
    assign S_out[71]  = A_iota[1][0][7];
    assign S_out[135]  = A_iota[2][0][7];
    assign S_out[199]  = A_iota[3][0][7];
    assign S_out[263]  = A_iota[4][0][7];
    assign S_out[327]  = A_iota[0][1][7];
    assign S_out[391]  = A_iota[1][1][7];
    assign S_out[455]  = A_iota[2][1][7];
    assign S_out[519]  = A_iota[3][1][7];
    assign S_out[583]  = A_iota[4][1][7];
    assign S_out[647]  = A_iota[0][2][7];
    assign S_out[711]  = A_iota[1][2][7];
    assign S_out[775]  = A_iota[2][2][7];
    assign S_out[839]  = A_iota[3][2][7];
    assign S_out[903]  = A_iota[4][2][7];
    assign S_out[967]  = A_iota[0][3][7];
    assign S_out[1031]  = A_iota[1][3][7];
    assign S_out[1095]  = A_iota[2][3][7];
    assign S_out[1159]  = A_iota[3][3][7];
    assign S_out[1223]  = A_iota[4][3][7];
    assign S_out[1287]  = A_iota[0][4][7];
    assign S_out[1351]  = A_iota[1][4][7];
    assign S_out[1415]  = A_iota[2][4][7];
    assign S_out[1479]  = A_iota[3][4][7];
    assign S_out[1543]  = A_iota[4][4][7];
    assign S_out[8]  = A_iota[0][0][8];
    assign S_out[72]  = A_iota[1][0][8];
    assign S_out[136]  = A_iota[2][0][8];
    assign S_out[200]  = A_iota[3][0][8];
    assign S_out[264]  = A_iota[4][0][8];
    assign S_out[328]  = A_iota[0][1][8];
    assign S_out[392]  = A_iota[1][1][8];
    assign S_out[456]  = A_iota[2][1][8];
    assign S_out[520]  = A_iota[3][1][8];
    assign S_out[584]  = A_iota[4][1][8];
    assign S_out[648]  = A_iota[0][2][8];
    assign S_out[712]  = A_iota[1][2][8];
    assign S_out[776]  = A_iota[2][2][8];
    assign S_out[840]  = A_iota[3][2][8];
    assign S_out[904]  = A_iota[4][2][8];
    assign S_out[968]  = A_iota[0][3][8];
    assign S_out[1032]  = A_iota[1][3][8];
    assign S_out[1096]  = A_iota[2][3][8];
    assign S_out[1160]  = A_iota[3][3][8];
    assign S_out[1224]  = A_iota[4][3][8];
    assign S_out[1288]  = A_iota[0][4][8];
    assign S_out[1352]  = A_iota[1][4][8];
    assign S_out[1416]  = A_iota[2][4][8];
    assign S_out[1480]  = A_iota[3][4][8];
    assign S_out[1544]  = A_iota[4][4][8];
    assign S_out[9]  = A_iota[0][0][9];
    assign S_out[73]  = A_iota[1][0][9];
    assign S_out[137]  = A_iota[2][0][9];
    assign S_out[201]  = A_iota[3][0][9];
    assign S_out[265]  = A_iota[4][0][9];
    assign S_out[329]  = A_iota[0][1][9];
    assign S_out[393]  = A_iota[1][1][9];
    assign S_out[457]  = A_iota[2][1][9];
    assign S_out[521]  = A_iota[3][1][9];
    assign S_out[585]  = A_iota[4][1][9];
    assign S_out[649]  = A_iota[0][2][9];
    assign S_out[713]  = A_iota[1][2][9];
    assign S_out[777]  = A_iota[2][2][9];
    assign S_out[841]  = A_iota[3][2][9];
    assign S_out[905]  = A_iota[4][2][9];
    assign S_out[969]  = A_iota[0][3][9];
    assign S_out[1033]  = A_iota[1][3][9];
    assign S_out[1097]  = A_iota[2][3][9];
    assign S_out[1161]  = A_iota[3][3][9];
    assign S_out[1225]  = A_iota[4][3][9];
    assign S_out[1289]  = A_iota[0][4][9];
    assign S_out[1353]  = A_iota[1][4][9];
    assign S_out[1417]  = A_iota[2][4][9];
    assign S_out[1481]  = A_iota[3][4][9];
    assign S_out[1545]  = A_iota[4][4][9];
    assign S_out[10]  = A_iota[0][0][10];
    assign S_out[74]  = A_iota[1][0][10];
    assign S_out[138]  = A_iota[2][0][10];
    assign S_out[202]  = A_iota[3][0][10];
    assign S_out[266]  = A_iota[4][0][10];
    assign S_out[330]  = A_iota[0][1][10];
    assign S_out[394]  = A_iota[1][1][10];
    assign S_out[458]  = A_iota[2][1][10];
    assign S_out[522]  = A_iota[3][1][10];
    assign S_out[586]  = A_iota[4][1][10];
    assign S_out[650]  = A_iota[0][2][10];
    assign S_out[714]  = A_iota[1][2][10];
    assign S_out[778]  = A_iota[2][2][10];
    assign S_out[842]  = A_iota[3][2][10];
    assign S_out[906]  = A_iota[4][2][10];
    assign S_out[970]  = A_iota[0][3][10];
    assign S_out[1034]  = A_iota[1][3][10];
    assign S_out[1098]  = A_iota[2][3][10];
    assign S_out[1162]  = A_iota[3][3][10];
    assign S_out[1226]  = A_iota[4][3][10];
    assign S_out[1290]  = A_iota[0][4][10];
    assign S_out[1354]  = A_iota[1][4][10];
    assign S_out[1418]  = A_iota[2][4][10];
    assign S_out[1482]  = A_iota[3][4][10];
    assign S_out[1546]  = A_iota[4][4][10];
    assign S_out[11]  = A_iota[0][0][11];
    assign S_out[75]  = A_iota[1][0][11];
    assign S_out[139]  = A_iota[2][0][11];
    assign S_out[203]  = A_iota[3][0][11];
    assign S_out[267]  = A_iota[4][0][11];
    assign S_out[331]  = A_iota[0][1][11];
    assign S_out[395]  = A_iota[1][1][11];
    assign S_out[459]  = A_iota[2][1][11];
    assign S_out[523]  = A_iota[3][1][11];
    assign S_out[587]  = A_iota[4][1][11];
    assign S_out[651]  = A_iota[0][2][11];
    assign S_out[715]  = A_iota[1][2][11];
    assign S_out[779]  = A_iota[2][2][11];
    assign S_out[843]  = A_iota[3][2][11];
    assign S_out[907]  = A_iota[4][2][11];
    assign S_out[971]  = A_iota[0][3][11];
    assign S_out[1035]  = A_iota[1][3][11];
    assign S_out[1099]  = A_iota[2][3][11];
    assign S_out[1163]  = A_iota[3][3][11];
    assign S_out[1227]  = A_iota[4][3][11];
    assign S_out[1291]  = A_iota[0][4][11];
    assign S_out[1355]  = A_iota[1][4][11];
    assign S_out[1419]  = A_iota[2][4][11];
    assign S_out[1483]  = A_iota[3][4][11];
    assign S_out[1547]  = A_iota[4][4][11];
    assign S_out[12]  = A_iota[0][0][12];
    assign S_out[76]  = A_iota[1][0][12];
    assign S_out[140]  = A_iota[2][0][12];
    assign S_out[204]  = A_iota[3][0][12];
    assign S_out[268]  = A_iota[4][0][12];
    assign S_out[332]  = A_iota[0][1][12];
    assign S_out[396]  = A_iota[1][1][12];
    assign S_out[460]  = A_iota[2][1][12];
    assign S_out[524]  = A_iota[3][1][12];
    assign S_out[588]  = A_iota[4][1][12];
    assign S_out[652]  = A_iota[0][2][12];
    assign S_out[716]  = A_iota[1][2][12];
    assign S_out[780]  = A_iota[2][2][12];
    assign S_out[844]  = A_iota[3][2][12];
    assign S_out[908]  = A_iota[4][2][12];
    assign S_out[972]  = A_iota[0][3][12];
    assign S_out[1036]  = A_iota[1][3][12];
    assign S_out[1100]  = A_iota[2][3][12];
    assign S_out[1164]  = A_iota[3][3][12];
    assign S_out[1228]  = A_iota[4][3][12];
    assign S_out[1292]  = A_iota[0][4][12];
    assign S_out[1356]  = A_iota[1][4][12];
    assign S_out[1420]  = A_iota[2][4][12];
    assign S_out[1484]  = A_iota[3][4][12];
    assign S_out[1548]  = A_iota[4][4][12];
    assign S_out[13]  = A_iota[0][0][13];
    assign S_out[77]  = A_iota[1][0][13];
    assign S_out[141]  = A_iota[2][0][13];
    assign S_out[205]  = A_iota[3][0][13];
    assign S_out[269]  = A_iota[4][0][13];
    assign S_out[333]  = A_iota[0][1][13];
    assign S_out[397]  = A_iota[1][1][13];
    assign S_out[461]  = A_iota[2][1][13];
    assign S_out[525]  = A_iota[3][1][13];
    assign S_out[589]  = A_iota[4][1][13];
    assign S_out[653]  = A_iota[0][2][13];
    assign S_out[717]  = A_iota[1][2][13];
    assign S_out[781]  = A_iota[2][2][13];
    assign S_out[845]  = A_iota[3][2][13];
    assign S_out[909]  = A_iota[4][2][13];
    assign S_out[973]  = A_iota[0][3][13];
    assign S_out[1037]  = A_iota[1][3][13];
    assign S_out[1101]  = A_iota[2][3][13];
    assign S_out[1165]  = A_iota[3][3][13];
    assign S_out[1229]  = A_iota[4][3][13];
    assign S_out[1293]  = A_iota[0][4][13];
    assign S_out[1357]  = A_iota[1][4][13];
    assign S_out[1421]  = A_iota[2][4][13];
    assign S_out[1485]  = A_iota[3][4][13];
    assign S_out[1549]  = A_iota[4][4][13];
    assign S_out[14]  = A_iota[0][0][14];
    assign S_out[78]  = A_iota[1][0][14];
    assign S_out[142]  = A_iota[2][0][14];
    assign S_out[206]  = A_iota[3][0][14];
    assign S_out[270]  = A_iota[4][0][14];
    assign S_out[334]  = A_iota[0][1][14];
    assign S_out[398]  = A_iota[1][1][14];
    assign S_out[462]  = A_iota[2][1][14];
    assign S_out[526]  = A_iota[3][1][14];
    assign S_out[590]  = A_iota[4][1][14];
    assign S_out[654]  = A_iota[0][2][14];
    assign S_out[718]  = A_iota[1][2][14];
    assign S_out[782]  = A_iota[2][2][14];
    assign S_out[846]  = A_iota[3][2][14];
    assign S_out[910]  = A_iota[4][2][14];
    assign S_out[974]  = A_iota[0][3][14];
    assign S_out[1038]  = A_iota[1][3][14];
    assign S_out[1102]  = A_iota[2][3][14];
    assign S_out[1166]  = A_iota[3][3][14];
    assign S_out[1230]  = A_iota[4][3][14];
    assign S_out[1294]  = A_iota[0][4][14];
    assign S_out[1358]  = A_iota[1][4][14];
    assign S_out[1422]  = A_iota[2][4][14];
    assign S_out[1486]  = A_iota[3][4][14];
    assign S_out[1550]  = A_iota[4][4][14];
    assign S_out[15]  = A_iota[0][0][15];
    assign S_out[79]  = A_iota[1][0][15];
    assign S_out[143]  = A_iota[2][0][15];
    assign S_out[207]  = A_iota[3][0][15];
    assign S_out[271]  = A_iota[4][0][15];
    assign S_out[335]  = A_iota[0][1][15];
    assign S_out[399]  = A_iota[1][1][15];
    assign S_out[463]  = A_iota[2][1][15];
    assign S_out[527]  = A_iota[3][1][15];
    assign S_out[591]  = A_iota[4][1][15];
    assign S_out[655]  = A_iota[0][2][15];
    assign S_out[719]  = A_iota[1][2][15];
    assign S_out[783]  = A_iota[2][2][15];
    assign S_out[847]  = A_iota[3][2][15];
    assign S_out[911]  = A_iota[4][2][15];
    assign S_out[975]  = A_iota[0][3][15];
    assign S_out[1039]  = A_iota[1][3][15];
    assign S_out[1103]  = A_iota[2][3][15];
    assign S_out[1167]  = A_iota[3][3][15];
    assign S_out[1231]  = A_iota[4][3][15];
    assign S_out[1295]  = A_iota[0][4][15];
    assign S_out[1359]  = A_iota[1][4][15];
    assign S_out[1423]  = A_iota[2][4][15];
    assign S_out[1487]  = A_iota[3][4][15];
    assign S_out[1551]  = A_iota[4][4][15];
    assign S_out[16]  = A_iota[0][0][16];
    assign S_out[80]  = A_iota[1][0][16];
    assign S_out[144]  = A_iota[2][0][16];
    assign S_out[208]  = A_iota[3][0][16];
    assign S_out[272]  = A_iota[4][0][16];
    assign S_out[336]  = A_iota[0][1][16];
    assign S_out[400]  = A_iota[1][1][16];
    assign S_out[464]  = A_iota[2][1][16];
    assign S_out[528]  = A_iota[3][1][16];
    assign S_out[592]  = A_iota[4][1][16];
    assign S_out[656]  = A_iota[0][2][16];
    assign S_out[720]  = A_iota[1][2][16];
    assign S_out[784]  = A_iota[2][2][16];
    assign S_out[848]  = A_iota[3][2][16];
    assign S_out[912]  = A_iota[4][2][16];
    assign S_out[976]  = A_iota[0][3][16];
    assign S_out[1040]  = A_iota[1][3][16];
    assign S_out[1104]  = A_iota[2][3][16];
    assign S_out[1168]  = A_iota[3][3][16];
    assign S_out[1232]  = A_iota[4][3][16];
    assign S_out[1296]  = A_iota[0][4][16];
    assign S_out[1360]  = A_iota[1][4][16];
    assign S_out[1424]  = A_iota[2][4][16];
    assign S_out[1488]  = A_iota[3][4][16];
    assign S_out[1552]  = A_iota[4][4][16];
    assign S_out[17]  = A_iota[0][0][17];
    assign S_out[81]  = A_iota[1][0][17];
    assign S_out[145]  = A_iota[2][0][17];
    assign S_out[209]  = A_iota[3][0][17];
    assign S_out[273]  = A_iota[4][0][17];
    assign S_out[337]  = A_iota[0][1][17];
    assign S_out[401]  = A_iota[1][1][17];
    assign S_out[465]  = A_iota[2][1][17];
    assign S_out[529]  = A_iota[3][1][17];
    assign S_out[593]  = A_iota[4][1][17];
    assign S_out[657]  = A_iota[0][2][17];
    assign S_out[721]  = A_iota[1][2][17];
    assign S_out[785]  = A_iota[2][2][17];
    assign S_out[849]  = A_iota[3][2][17];
    assign S_out[913]  = A_iota[4][2][17];
    assign S_out[977]  = A_iota[0][3][17];
    assign S_out[1041]  = A_iota[1][3][17];
    assign S_out[1105]  = A_iota[2][3][17];
    assign S_out[1169]  = A_iota[3][3][17];
    assign S_out[1233]  = A_iota[4][3][17];
    assign S_out[1297]  = A_iota[0][4][17];
    assign S_out[1361]  = A_iota[1][4][17];
    assign S_out[1425]  = A_iota[2][4][17];
    assign S_out[1489]  = A_iota[3][4][17];
    assign S_out[1553]  = A_iota[4][4][17];
    assign S_out[18]  = A_iota[0][0][18];
    assign S_out[82]  = A_iota[1][0][18];
    assign S_out[146]  = A_iota[2][0][18];
    assign S_out[210]  = A_iota[3][0][18];
    assign S_out[274]  = A_iota[4][0][18];
    assign S_out[338]  = A_iota[0][1][18];
    assign S_out[402]  = A_iota[1][1][18];
    assign S_out[466]  = A_iota[2][1][18];
    assign S_out[530]  = A_iota[3][1][18];
    assign S_out[594]  = A_iota[4][1][18];
    assign S_out[658]  = A_iota[0][2][18];
    assign S_out[722]  = A_iota[1][2][18];
    assign S_out[786]  = A_iota[2][2][18];
    assign S_out[850]  = A_iota[3][2][18];
    assign S_out[914]  = A_iota[4][2][18];
    assign S_out[978]  = A_iota[0][3][18];
    assign S_out[1042]  = A_iota[1][3][18];
    assign S_out[1106]  = A_iota[2][3][18];
    assign S_out[1170]  = A_iota[3][3][18];
    assign S_out[1234]  = A_iota[4][3][18];
    assign S_out[1298]  = A_iota[0][4][18];
    assign S_out[1362]  = A_iota[1][4][18];
    assign S_out[1426]  = A_iota[2][4][18];
    assign S_out[1490]  = A_iota[3][4][18];
    assign S_out[1554]  = A_iota[4][4][18];
    assign S_out[19]  = A_iota[0][0][19];
    assign S_out[83]  = A_iota[1][0][19];
    assign S_out[147]  = A_iota[2][0][19];
    assign S_out[211]  = A_iota[3][0][19];
    assign S_out[275]  = A_iota[4][0][19];
    assign S_out[339]  = A_iota[0][1][19];
    assign S_out[403]  = A_iota[1][1][19];
    assign S_out[467]  = A_iota[2][1][19];
    assign S_out[531]  = A_iota[3][1][19];
    assign S_out[595]  = A_iota[4][1][19];
    assign S_out[659]  = A_iota[0][2][19];
    assign S_out[723]  = A_iota[1][2][19];
    assign S_out[787]  = A_iota[2][2][19];
    assign S_out[851]  = A_iota[3][2][19];
    assign S_out[915]  = A_iota[4][2][19];
    assign S_out[979]  = A_iota[0][3][19];
    assign S_out[1043]  = A_iota[1][3][19];
    assign S_out[1107]  = A_iota[2][3][19];
    assign S_out[1171]  = A_iota[3][3][19];
    assign S_out[1235]  = A_iota[4][3][19];
    assign S_out[1299]  = A_iota[0][4][19];
    assign S_out[1363]  = A_iota[1][4][19];
    assign S_out[1427]  = A_iota[2][4][19];
    assign S_out[1491]  = A_iota[3][4][19];
    assign S_out[1555]  = A_iota[4][4][19];
    assign S_out[20]  = A_iota[0][0][20];
    assign S_out[84]  = A_iota[1][0][20];
    assign S_out[148]  = A_iota[2][0][20];
    assign S_out[212]  = A_iota[3][0][20];
    assign S_out[276]  = A_iota[4][0][20];
    assign S_out[340]  = A_iota[0][1][20];
    assign S_out[404]  = A_iota[1][1][20];
    assign S_out[468]  = A_iota[2][1][20];
    assign S_out[532]  = A_iota[3][1][20];
    assign S_out[596]  = A_iota[4][1][20];
    assign S_out[660]  = A_iota[0][2][20];
    assign S_out[724]  = A_iota[1][2][20];
    assign S_out[788]  = A_iota[2][2][20];
    assign S_out[852]  = A_iota[3][2][20];
    assign S_out[916]  = A_iota[4][2][20];
    assign S_out[980]  = A_iota[0][3][20];
    assign S_out[1044]  = A_iota[1][3][20];
    assign S_out[1108]  = A_iota[2][3][20];
    assign S_out[1172]  = A_iota[3][3][20];
    assign S_out[1236]  = A_iota[4][3][20];
    assign S_out[1300]  = A_iota[0][4][20];
    assign S_out[1364]  = A_iota[1][4][20];
    assign S_out[1428]  = A_iota[2][4][20];
    assign S_out[1492]  = A_iota[3][4][20];
    assign S_out[1556]  = A_iota[4][4][20];
    assign S_out[21]  = A_iota[0][0][21];
    assign S_out[85]  = A_iota[1][0][21];
    assign S_out[149]  = A_iota[2][0][21];
    assign S_out[213]  = A_iota[3][0][21];
    assign S_out[277]  = A_iota[4][0][21];
    assign S_out[341]  = A_iota[0][1][21];
    assign S_out[405]  = A_iota[1][1][21];
    assign S_out[469]  = A_iota[2][1][21];
    assign S_out[533]  = A_iota[3][1][21];
    assign S_out[597]  = A_iota[4][1][21];
    assign S_out[661]  = A_iota[0][2][21];
    assign S_out[725]  = A_iota[1][2][21];
    assign S_out[789]  = A_iota[2][2][21];
    assign S_out[853]  = A_iota[3][2][21];
    assign S_out[917]  = A_iota[4][2][21];
    assign S_out[981]  = A_iota[0][3][21];
    assign S_out[1045]  = A_iota[1][3][21];
    assign S_out[1109]  = A_iota[2][3][21];
    assign S_out[1173]  = A_iota[3][3][21];
    assign S_out[1237]  = A_iota[4][3][21];
    assign S_out[1301]  = A_iota[0][4][21];
    assign S_out[1365]  = A_iota[1][4][21];
    assign S_out[1429]  = A_iota[2][4][21];
    assign S_out[1493]  = A_iota[3][4][21];
    assign S_out[1557]  = A_iota[4][4][21];
    assign S_out[22]  = A_iota[0][0][22];
    assign S_out[86]  = A_iota[1][0][22];
    assign S_out[150]  = A_iota[2][0][22];
    assign S_out[214]  = A_iota[3][0][22];
    assign S_out[278]  = A_iota[4][0][22];
    assign S_out[342]  = A_iota[0][1][22];
    assign S_out[406]  = A_iota[1][1][22];
    assign S_out[470]  = A_iota[2][1][22];
    assign S_out[534]  = A_iota[3][1][22];
    assign S_out[598]  = A_iota[4][1][22];
    assign S_out[662]  = A_iota[0][2][22];
    assign S_out[726]  = A_iota[1][2][22];
    assign S_out[790]  = A_iota[2][2][22];
    assign S_out[854]  = A_iota[3][2][22];
    assign S_out[918]  = A_iota[4][2][22];
    assign S_out[982]  = A_iota[0][3][22];
    assign S_out[1046]  = A_iota[1][3][22];
    assign S_out[1110]  = A_iota[2][3][22];
    assign S_out[1174]  = A_iota[3][3][22];
    assign S_out[1238]  = A_iota[4][3][22];
    assign S_out[1302]  = A_iota[0][4][22];
    assign S_out[1366]  = A_iota[1][4][22];
    assign S_out[1430]  = A_iota[2][4][22];
    assign S_out[1494]  = A_iota[3][4][22];
    assign S_out[1558]  = A_iota[4][4][22];
    assign S_out[23]  = A_iota[0][0][23];
    assign S_out[87]  = A_iota[1][0][23];
    assign S_out[151]  = A_iota[2][0][23];
    assign S_out[215]  = A_iota[3][0][23];
    assign S_out[279]  = A_iota[4][0][23];
    assign S_out[343]  = A_iota[0][1][23];
    assign S_out[407]  = A_iota[1][1][23];
    assign S_out[471]  = A_iota[2][1][23];
    assign S_out[535]  = A_iota[3][1][23];
    assign S_out[599]  = A_iota[4][1][23];
    assign S_out[663]  = A_iota[0][2][23];
    assign S_out[727]  = A_iota[1][2][23];
    assign S_out[791]  = A_iota[2][2][23];
    assign S_out[855]  = A_iota[3][2][23];
    assign S_out[919]  = A_iota[4][2][23];
    assign S_out[983]  = A_iota[0][3][23];
    assign S_out[1047]  = A_iota[1][3][23];
    assign S_out[1111]  = A_iota[2][3][23];
    assign S_out[1175]  = A_iota[3][3][23];
    assign S_out[1239]  = A_iota[4][3][23];
    assign S_out[1303]  = A_iota[0][4][23];
    assign S_out[1367]  = A_iota[1][4][23];
    assign S_out[1431]  = A_iota[2][4][23];
    assign S_out[1495]  = A_iota[3][4][23];
    assign S_out[1559]  = A_iota[4][4][23];
    assign S_out[24]  = A_iota[0][0][24];
    assign S_out[88]  = A_iota[1][0][24];
    assign S_out[152]  = A_iota[2][0][24];
    assign S_out[216]  = A_iota[3][0][24];
    assign S_out[280]  = A_iota[4][0][24];
    assign S_out[344]  = A_iota[0][1][24];
    assign S_out[408]  = A_iota[1][1][24];
    assign S_out[472]  = A_iota[2][1][24];
    assign S_out[536]  = A_iota[3][1][24];
    assign S_out[600]  = A_iota[4][1][24];
    assign S_out[664]  = A_iota[0][2][24];
    assign S_out[728]  = A_iota[1][2][24];
    assign S_out[792]  = A_iota[2][2][24];
    assign S_out[856]  = A_iota[3][2][24];
    assign S_out[920]  = A_iota[4][2][24];
    assign S_out[984]  = A_iota[0][3][24];
    assign S_out[1048]  = A_iota[1][3][24];
    assign S_out[1112]  = A_iota[2][3][24];
    assign S_out[1176]  = A_iota[3][3][24];
    assign S_out[1240]  = A_iota[4][3][24];
    assign S_out[1304]  = A_iota[0][4][24];
    assign S_out[1368]  = A_iota[1][4][24];
    assign S_out[1432]  = A_iota[2][4][24];
    assign S_out[1496]  = A_iota[3][4][24];
    assign S_out[1560]  = A_iota[4][4][24];
    assign S_out[25]  = A_iota[0][0][25];
    assign S_out[89]  = A_iota[1][0][25];
    assign S_out[153]  = A_iota[2][0][25];
    assign S_out[217]  = A_iota[3][0][25];
    assign S_out[281]  = A_iota[4][0][25];
    assign S_out[345]  = A_iota[0][1][25];
    assign S_out[409]  = A_iota[1][1][25];
    assign S_out[473]  = A_iota[2][1][25];
    assign S_out[537]  = A_iota[3][1][25];
    assign S_out[601]  = A_iota[4][1][25];
    assign S_out[665]  = A_iota[0][2][25];
    assign S_out[729]  = A_iota[1][2][25];
    assign S_out[793]  = A_iota[2][2][25];
    assign S_out[857]  = A_iota[3][2][25];
    assign S_out[921]  = A_iota[4][2][25];
    assign S_out[985]  = A_iota[0][3][25];
    assign S_out[1049]  = A_iota[1][3][25];
    assign S_out[1113]  = A_iota[2][3][25];
    assign S_out[1177]  = A_iota[3][3][25];
    assign S_out[1241]  = A_iota[4][3][25];
    assign S_out[1305]  = A_iota[0][4][25];
    assign S_out[1369]  = A_iota[1][4][25];
    assign S_out[1433]  = A_iota[2][4][25];
    assign S_out[1497]  = A_iota[3][4][25];
    assign S_out[1561]  = A_iota[4][4][25];
    assign S_out[26]  = A_iota[0][0][26];
    assign S_out[90]  = A_iota[1][0][26];
    assign S_out[154]  = A_iota[2][0][26];
    assign S_out[218]  = A_iota[3][0][26];
    assign S_out[282]  = A_iota[4][0][26];
    assign S_out[346]  = A_iota[0][1][26];
    assign S_out[410]  = A_iota[1][1][26];
    assign S_out[474]  = A_iota[2][1][26];
    assign S_out[538]  = A_iota[3][1][26];
    assign S_out[602]  = A_iota[4][1][26];
    assign S_out[666]  = A_iota[0][2][26];
    assign S_out[730]  = A_iota[1][2][26];
    assign S_out[794]  = A_iota[2][2][26];
    assign S_out[858]  = A_iota[3][2][26];
    assign S_out[922]  = A_iota[4][2][26];
    assign S_out[986]  = A_iota[0][3][26];
    assign S_out[1050]  = A_iota[1][3][26];
    assign S_out[1114]  = A_iota[2][3][26];
    assign S_out[1178]  = A_iota[3][3][26];
    assign S_out[1242]  = A_iota[4][3][26];
    assign S_out[1306]  = A_iota[0][4][26];
    assign S_out[1370]  = A_iota[1][4][26];
    assign S_out[1434]  = A_iota[2][4][26];
    assign S_out[1498]  = A_iota[3][4][26];
    assign S_out[1562]  = A_iota[4][4][26];
    assign S_out[27]  = A_iota[0][0][27];
    assign S_out[91]  = A_iota[1][0][27];
    assign S_out[155]  = A_iota[2][0][27];
    assign S_out[219]  = A_iota[3][0][27];
    assign S_out[283]  = A_iota[4][0][27];
    assign S_out[347]  = A_iota[0][1][27];
    assign S_out[411]  = A_iota[1][1][27];
    assign S_out[475]  = A_iota[2][1][27];
    assign S_out[539]  = A_iota[3][1][27];
    assign S_out[603]  = A_iota[4][1][27];
    assign S_out[667]  = A_iota[0][2][27];
    assign S_out[731]  = A_iota[1][2][27];
    assign S_out[795]  = A_iota[2][2][27];
    assign S_out[859]  = A_iota[3][2][27];
    assign S_out[923]  = A_iota[4][2][27];
    assign S_out[987]  = A_iota[0][3][27];
    assign S_out[1051]  = A_iota[1][3][27];
    assign S_out[1115]  = A_iota[2][3][27];
    assign S_out[1179]  = A_iota[3][3][27];
    assign S_out[1243]  = A_iota[4][3][27];
    assign S_out[1307]  = A_iota[0][4][27];
    assign S_out[1371]  = A_iota[1][4][27];
    assign S_out[1435]  = A_iota[2][4][27];
    assign S_out[1499]  = A_iota[3][4][27];
    assign S_out[1563]  = A_iota[4][4][27];
    assign S_out[28]  = A_iota[0][0][28];
    assign S_out[92]  = A_iota[1][0][28];
    assign S_out[156]  = A_iota[2][0][28];
    assign S_out[220]  = A_iota[3][0][28];
    assign S_out[284]  = A_iota[4][0][28];
    assign S_out[348]  = A_iota[0][1][28];
    assign S_out[412]  = A_iota[1][1][28];
    assign S_out[476]  = A_iota[2][1][28];
    assign S_out[540]  = A_iota[3][1][28];
    assign S_out[604]  = A_iota[4][1][28];
    assign S_out[668]  = A_iota[0][2][28];
    assign S_out[732]  = A_iota[1][2][28];
    assign S_out[796]  = A_iota[2][2][28];
    assign S_out[860]  = A_iota[3][2][28];
    assign S_out[924]  = A_iota[4][2][28];
    assign S_out[988]  = A_iota[0][3][28];
    assign S_out[1052]  = A_iota[1][3][28];
    assign S_out[1116]  = A_iota[2][3][28];
    assign S_out[1180]  = A_iota[3][3][28];
    assign S_out[1244]  = A_iota[4][3][28];
    assign S_out[1308]  = A_iota[0][4][28];
    assign S_out[1372]  = A_iota[1][4][28];
    assign S_out[1436]  = A_iota[2][4][28];
    assign S_out[1500]  = A_iota[3][4][28];
    assign S_out[1564]  = A_iota[4][4][28];
    assign S_out[29]  = A_iota[0][0][29];
    assign S_out[93]  = A_iota[1][0][29];
    assign S_out[157]  = A_iota[2][0][29];
    assign S_out[221]  = A_iota[3][0][29];
    assign S_out[285]  = A_iota[4][0][29];
    assign S_out[349]  = A_iota[0][1][29];
    assign S_out[413]  = A_iota[1][1][29];
    assign S_out[477]  = A_iota[2][1][29];
    assign S_out[541]  = A_iota[3][1][29];
    assign S_out[605]  = A_iota[4][1][29];
    assign S_out[669]  = A_iota[0][2][29];
    assign S_out[733]  = A_iota[1][2][29];
    assign S_out[797]  = A_iota[2][2][29];
    assign S_out[861]  = A_iota[3][2][29];
    assign S_out[925]  = A_iota[4][2][29];
    assign S_out[989]  = A_iota[0][3][29];
    assign S_out[1053]  = A_iota[1][3][29];
    assign S_out[1117]  = A_iota[2][3][29];
    assign S_out[1181]  = A_iota[3][3][29];
    assign S_out[1245]  = A_iota[4][3][29];
    assign S_out[1309]  = A_iota[0][4][29];
    assign S_out[1373]  = A_iota[1][4][29];
    assign S_out[1437]  = A_iota[2][4][29];
    assign S_out[1501]  = A_iota[3][4][29];
    assign S_out[1565]  = A_iota[4][4][29];
    assign S_out[30]  = A_iota[0][0][30];
    assign S_out[94]  = A_iota[1][0][30];
    assign S_out[158]  = A_iota[2][0][30];
    assign S_out[222]  = A_iota[3][0][30];
    assign S_out[286]  = A_iota[4][0][30];
    assign S_out[350]  = A_iota[0][1][30];
    assign S_out[414]  = A_iota[1][1][30];
    assign S_out[478]  = A_iota[2][1][30];
    assign S_out[542]  = A_iota[3][1][30];
    assign S_out[606]  = A_iota[4][1][30];
    assign S_out[670]  = A_iota[0][2][30];
    assign S_out[734]  = A_iota[1][2][30];
    assign S_out[798]  = A_iota[2][2][30];
    assign S_out[862]  = A_iota[3][2][30];
    assign S_out[926]  = A_iota[4][2][30];
    assign S_out[990]  = A_iota[0][3][30];
    assign S_out[1054]  = A_iota[1][3][30];
    assign S_out[1118]  = A_iota[2][3][30];
    assign S_out[1182]  = A_iota[3][3][30];
    assign S_out[1246]  = A_iota[4][3][30];
    assign S_out[1310]  = A_iota[0][4][30];
    assign S_out[1374]  = A_iota[1][4][30];
    assign S_out[1438]  = A_iota[2][4][30];
    assign S_out[1502]  = A_iota[3][4][30];
    assign S_out[1566]  = A_iota[4][4][30];
    assign S_out[31]  = A_iota[0][0][31];
    assign S_out[95]  = A_iota[1][0][31];
    assign S_out[159]  = A_iota[2][0][31];
    assign S_out[223]  = A_iota[3][0][31];
    assign S_out[287]  = A_iota[4][0][31];
    assign S_out[351]  = A_iota[0][1][31];
    assign S_out[415]  = A_iota[1][1][31];
    assign S_out[479]  = A_iota[2][1][31];
    assign S_out[543]  = A_iota[3][1][31];
    assign S_out[607]  = A_iota[4][1][31];
    assign S_out[671]  = A_iota[0][2][31];
    assign S_out[735]  = A_iota[1][2][31];
    assign S_out[799]  = A_iota[2][2][31];
    assign S_out[863]  = A_iota[3][2][31];
    assign S_out[927]  = A_iota[4][2][31];
    assign S_out[991]  = A_iota[0][3][31];
    assign S_out[1055]  = A_iota[1][3][31];
    assign S_out[1119]  = A_iota[2][3][31];
    assign S_out[1183]  = A_iota[3][3][31];
    assign S_out[1247]  = A_iota[4][3][31];
    assign S_out[1311]  = A_iota[0][4][31];
    assign S_out[1375]  = A_iota[1][4][31];
    assign S_out[1439]  = A_iota[2][4][31];
    assign S_out[1503]  = A_iota[3][4][31];
    assign S_out[1567]  = A_iota[4][4][31];
    assign S_out[32]  = A_iota[0][0][32];
    assign S_out[96]  = A_iota[1][0][32];
    assign S_out[160]  = A_iota[2][0][32];
    assign S_out[224]  = A_iota[3][0][32];
    assign S_out[288]  = A_iota[4][0][32];
    assign S_out[352]  = A_iota[0][1][32];
    assign S_out[416]  = A_iota[1][1][32];
    assign S_out[480]  = A_iota[2][1][32];
    assign S_out[544]  = A_iota[3][1][32];
    assign S_out[608]  = A_iota[4][1][32];
    assign S_out[672]  = A_iota[0][2][32];
    assign S_out[736]  = A_iota[1][2][32];
    assign S_out[800]  = A_iota[2][2][32];
    assign S_out[864]  = A_iota[3][2][32];
    assign S_out[928]  = A_iota[4][2][32];
    assign S_out[992]  = A_iota[0][3][32];
    assign S_out[1056]  = A_iota[1][3][32];
    assign S_out[1120]  = A_iota[2][3][32];
    assign S_out[1184]  = A_iota[3][3][32];
    assign S_out[1248]  = A_iota[4][3][32];
    assign S_out[1312]  = A_iota[0][4][32];
    assign S_out[1376]  = A_iota[1][4][32];
    assign S_out[1440]  = A_iota[2][4][32];
    assign S_out[1504]  = A_iota[3][4][32];
    assign S_out[1568]  = A_iota[4][4][32];
    assign S_out[33]  = A_iota[0][0][33];
    assign S_out[97]  = A_iota[1][0][33];
    assign S_out[161]  = A_iota[2][0][33];
    assign S_out[225]  = A_iota[3][0][33];
    assign S_out[289]  = A_iota[4][0][33];
    assign S_out[353]  = A_iota[0][1][33];
    assign S_out[417]  = A_iota[1][1][33];
    assign S_out[481]  = A_iota[2][1][33];
    assign S_out[545]  = A_iota[3][1][33];
    assign S_out[609]  = A_iota[4][1][33];
    assign S_out[673]  = A_iota[0][2][33];
    assign S_out[737]  = A_iota[1][2][33];
    assign S_out[801]  = A_iota[2][2][33];
    assign S_out[865]  = A_iota[3][2][33];
    assign S_out[929]  = A_iota[4][2][33];
    assign S_out[993]  = A_iota[0][3][33];
    assign S_out[1057]  = A_iota[1][3][33];
    assign S_out[1121]  = A_iota[2][3][33];
    assign S_out[1185]  = A_iota[3][3][33];
    assign S_out[1249]  = A_iota[4][3][33];
    assign S_out[1313]  = A_iota[0][4][33];
    assign S_out[1377]  = A_iota[1][4][33];
    assign S_out[1441]  = A_iota[2][4][33];
    assign S_out[1505]  = A_iota[3][4][33];
    assign S_out[1569]  = A_iota[4][4][33];
    assign S_out[34]  = A_iota[0][0][34];
    assign S_out[98]  = A_iota[1][0][34];
    assign S_out[162]  = A_iota[2][0][34];
    assign S_out[226]  = A_iota[3][0][34];
    assign S_out[290]  = A_iota[4][0][34];
    assign S_out[354]  = A_iota[0][1][34];
    assign S_out[418]  = A_iota[1][1][34];
    assign S_out[482]  = A_iota[2][1][34];
    assign S_out[546]  = A_iota[3][1][34];
    assign S_out[610]  = A_iota[4][1][34];
    assign S_out[674]  = A_iota[0][2][34];
    assign S_out[738]  = A_iota[1][2][34];
    assign S_out[802]  = A_iota[2][2][34];
    assign S_out[866]  = A_iota[3][2][34];
    assign S_out[930]  = A_iota[4][2][34];
    assign S_out[994]  = A_iota[0][3][34];
    assign S_out[1058]  = A_iota[1][3][34];
    assign S_out[1122]  = A_iota[2][3][34];
    assign S_out[1186]  = A_iota[3][3][34];
    assign S_out[1250]  = A_iota[4][3][34];
    assign S_out[1314]  = A_iota[0][4][34];
    assign S_out[1378]  = A_iota[1][4][34];
    assign S_out[1442]  = A_iota[2][4][34];
    assign S_out[1506]  = A_iota[3][4][34];
    assign S_out[1570]  = A_iota[4][4][34];
    assign S_out[35]  = A_iota[0][0][35];
    assign S_out[99]  = A_iota[1][0][35];
    assign S_out[163]  = A_iota[2][0][35];
    assign S_out[227]  = A_iota[3][0][35];
    assign S_out[291]  = A_iota[4][0][35];
    assign S_out[355]  = A_iota[0][1][35];
    assign S_out[419]  = A_iota[1][1][35];
    assign S_out[483]  = A_iota[2][1][35];
    assign S_out[547]  = A_iota[3][1][35];
    assign S_out[611]  = A_iota[4][1][35];
    assign S_out[675]  = A_iota[0][2][35];
    assign S_out[739]  = A_iota[1][2][35];
    assign S_out[803]  = A_iota[2][2][35];
    assign S_out[867]  = A_iota[3][2][35];
    assign S_out[931]  = A_iota[4][2][35];
    assign S_out[995]  = A_iota[0][3][35];
    assign S_out[1059]  = A_iota[1][3][35];
    assign S_out[1123]  = A_iota[2][3][35];
    assign S_out[1187]  = A_iota[3][3][35];
    assign S_out[1251]  = A_iota[4][3][35];
    assign S_out[1315]  = A_iota[0][4][35];
    assign S_out[1379]  = A_iota[1][4][35];
    assign S_out[1443]  = A_iota[2][4][35];
    assign S_out[1507]  = A_iota[3][4][35];
    assign S_out[1571]  = A_iota[4][4][35];
    assign S_out[36]  = A_iota[0][0][36];
    assign S_out[100]  = A_iota[1][0][36];
    assign S_out[164]  = A_iota[2][0][36];
    assign S_out[228]  = A_iota[3][0][36];
    assign S_out[292]  = A_iota[4][0][36];
    assign S_out[356]  = A_iota[0][1][36];
    assign S_out[420]  = A_iota[1][1][36];
    assign S_out[484]  = A_iota[2][1][36];
    assign S_out[548]  = A_iota[3][1][36];
    assign S_out[612]  = A_iota[4][1][36];
    assign S_out[676]  = A_iota[0][2][36];
    assign S_out[740]  = A_iota[1][2][36];
    assign S_out[804]  = A_iota[2][2][36];
    assign S_out[868]  = A_iota[3][2][36];
    assign S_out[932]  = A_iota[4][2][36];
    assign S_out[996]  = A_iota[0][3][36];
    assign S_out[1060]  = A_iota[1][3][36];
    assign S_out[1124]  = A_iota[2][3][36];
    assign S_out[1188]  = A_iota[3][3][36];
    assign S_out[1252]  = A_iota[4][3][36];
    assign S_out[1316]  = A_iota[0][4][36];
    assign S_out[1380]  = A_iota[1][4][36];
    assign S_out[1444]  = A_iota[2][4][36];
    assign S_out[1508]  = A_iota[3][4][36];
    assign S_out[1572]  = A_iota[4][4][36];
    assign S_out[37]  = A_iota[0][0][37];
    assign S_out[101]  = A_iota[1][0][37];
    assign S_out[165]  = A_iota[2][0][37];
    assign S_out[229]  = A_iota[3][0][37];
    assign S_out[293]  = A_iota[4][0][37];
    assign S_out[357]  = A_iota[0][1][37];
    assign S_out[421]  = A_iota[1][1][37];
    assign S_out[485]  = A_iota[2][1][37];
    assign S_out[549]  = A_iota[3][1][37];
    assign S_out[613]  = A_iota[4][1][37];
    assign S_out[677]  = A_iota[0][2][37];
    assign S_out[741]  = A_iota[1][2][37];
    assign S_out[805]  = A_iota[2][2][37];
    assign S_out[869]  = A_iota[3][2][37];
    assign S_out[933]  = A_iota[4][2][37];
    assign S_out[997]  = A_iota[0][3][37];
    assign S_out[1061]  = A_iota[1][3][37];
    assign S_out[1125]  = A_iota[2][3][37];
    assign S_out[1189]  = A_iota[3][3][37];
    assign S_out[1253]  = A_iota[4][3][37];
    assign S_out[1317]  = A_iota[0][4][37];
    assign S_out[1381]  = A_iota[1][4][37];
    assign S_out[1445]  = A_iota[2][4][37];
    assign S_out[1509]  = A_iota[3][4][37];
    assign S_out[1573]  = A_iota[4][4][37];
    assign S_out[38]  = A_iota[0][0][38];
    assign S_out[102]  = A_iota[1][0][38];
    assign S_out[166]  = A_iota[2][0][38];
    assign S_out[230]  = A_iota[3][0][38];
    assign S_out[294]  = A_iota[4][0][38];
    assign S_out[358]  = A_iota[0][1][38];
    assign S_out[422]  = A_iota[1][1][38];
    assign S_out[486]  = A_iota[2][1][38];
    assign S_out[550]  = A_iota[3][1][38];
    assign S_out[614]  = A_iota[4][1][38];
    assign S_out[678]  = A_iota[0][2][38];
    assign S_out[742]  = A_iota[1][2][38];
    assign S_out[806]  = A_iota[2][2][38];
    assign S_out[870]  = A_iota[3][2][38];
    assign S_out[934]  = A_iota[4][2][38];
    assign S_out[998]  = A_iota[0][3][38];
    assign S_out[1062]  = A_iota[1][3][38];
    assign S_out[1126]  = A_iota[2][3][38];
    assign S_out[1190]  = A_iota[3][3][38];
    assign S_out[1254]  = A_iota[4][3][38];
    assign S_out[1318]  = A_iota[0][4][38];
    assign S_out[1382]  = A_iota[1][4][38];
    assign S_out[1446]  = A_iota[2][4][38];
    assign S_out[1510]  = A_iota[3][4][38];
    assign S_out[1574]  = A_iota[4][4][38];
    assign S_out[39]  = A_iota[0][0][39];
    assign S_out[103]  = A_iota[1][0][39];
    assign S_out[167]  = A_iota[2][0][39];
    assign S_out[231]  = A_iota[3][0][39];
    assign S_out[295]  = A_iota[4][0][39];
    assign S_out[359]  = A_iota[0][1][39];
    assign S_out[423]  = A_iota[1][1][39];
    assign S_out[487]  = A_iota[2][1][39];
    assign S_out[551]  = A_iota[3][1][39];
    assign S_out[615]  = A_iota[4][1][39];
    assign S_out[679]  = A_iota[0][2][39];
    assign S_out[743]  = A_iota[1][2][39];
    assign S_out[807]  = A_iota[2][2][39];
    assign S_out[871]  = A_iota[3][2][39];
    assign S_out[935]  = A_iota[4][2][39];
    assign S_out[999]  = A_iota[0][3][39];
    assign S_out[1063]  = A_iota[1][3][39];
    assign S_out[1127]  = A_iota[2][3][39];
    assign S_out[1191]  = A_iota[3][3][39];
    assign S_out[1255]  = A_iota[4][3][39];
    assign S_out[1319]  = A_iota[0][4][39];
    assign S_out[1383]  = A_iota[1][4][39];
    assign S_out[1447]  = A_iota[2][4][39];
    assign S_out[1511]  = A_iota[3][4][39];
    assign S_out[1575]  = A_iota[4][4][39];
    assign S_out[40]  = A_iota[0][0][40];
    assign S_out[104]  = A_iota[1][0][40];
    assign S_out[168]  = A_iota[2][0][40];
    assign S_out[232]  = A_iota[3][0][40];
    assign S_out[296]  = A_iota[4][0][40];
    assign S_out[360]  = A_iota[0][1][40];
    assign S_out[424]  = A_iota[1][1][40];
    assign S_out[488]  = A_iota[2][1][40];
    assign S_out[552]  = A_iota[3][1][40];
    assign S_out[616]  = A_iota[4][1][40];
    assign S_out[680]  = A_iota[0][2][40];
    assign S_out[744]  = A_iota[1][2][40];
    assign S_out[808]  = A_iota[2][2][40];
    assign S_out[872]  = A_iota[3][2][40];
    assign S_out[936]  = A_iota[4][2][40];
    assign S_out[1000]  = A_iota[0][3][40];
    assign S_out[1064]  = A_iota[1][3][40];
    assign S_out[1128]  = A_iota[2][3][40];
    assign S_out[1192]  = A_iota[3][3][40];
    assign S_out[1256]  = A_iota[4][3][40];
    assign S_out[1320]  = A_iota[0][4][40];
    assign S_out[1384]  = A_iota[1][4][40];
    assign S_out[1448]  = A_iota[2][4][40];
    assign S_out[1512]  = A_iota[3][4][40];
    assign S_out[1576]  = A_iota[4][4][40];
    assign S_out[41]  = A_iota[0][0][41];
    assign S_out[105]  = A_iota[1][0][41];
    assign S_out[169]  = A_iota[2][0][41];
    assign S_out[233]  = A_iota[3][0][41];
    assign S_out[297]  = A_iota[4][0][41];
    assign S_out[361]  = A_iota[0][1][41];
    assign S_out[425]  = A_iota[1][1][41];
    assign S_out[489]  = A_iota[2][1][41];
    assign S_out[553]  = A_iota[3][1][41];
    assign S_out[617]  = A_iota[4][1][41];
    assign S_out[681]  = A_iota[0][2][41];
    assign S_out[745]  = A_iota[1][2][41];
    assign S_out[809]  = A_iota[2][2][41];
    assign S_out[873]  = A_iota[3][2][41];
    assign S_out[937]  = A_iota[4][2][41];
    assign S_out[1001]  = A_iota[0][3][41];
    assign S_out[1065]  = A_iota[1][3][41];
    assign S_out[1129]  = A_iota[2][3][41];
    assign S_out[1193]  = A_iota[3][3][41];
    assign S_out[1257]  = A_iota[4][3][41];
    assign S_out[1321]  = A_iota[0][4][41];
    assign S_out[1385]  = A_iota[1][4][41];
    assign S_out[1449]  = A_iota[2][4][41];
    assign S_out[1513]  = A_iota[3][4][41];
    assign S_out[1577]  = A_iota[4][4][41];
    assign S_out[42]  = A_iota[0][0][42];
    assign S_out[106]  = A_iota[1][0][42];
    assign S_out[170]  = A_iota[2][0][42];
    assign S_out[234]  = A_iota[3][0][42];
    assign S_out[298]  = A_iota[4][0][42];
    assign S_out[362]  = A_iota[0][1][42];
    assign S_out[426]  = A_iota[1][1][42];
    assign S_out[490]  = A_iota[2][1][42];
    assign S_out[554]  = A_iota[3][1][42];
    assign S_out[618]  = A_iota[4][1][42];
    assign S_out[682]  = A_iota[0][2][42];
    assign S_out[746]  = A_iota[1][2][42];
    assign S_out[810]  = A_iota[2][2][42];
    assign S_out[874]  = A_iota[3][2][42];
    assign S_out[938]  = A_iota[4][2][42];
    assign S_out[1002]  = A_iota[0][3][42];
    assign S_out[1066]  = A_iota[1][3][42];
    assign S_out[1130]  = A_iota[2][3][42];
    assign S_out[1194]  = A_iota[3][3][42];
    assign S_out[1258]  = A_iota[4][3][42];
    assign S_out[1322]  = A_iota[0][4][42];
    assign S_out[1386]  = A_iota[1][4][42];
    assign S_out[1450]  = A_iota[2][4][42];
    assign S_out[1514]  = A_iota[3][4][42];
    assign S_out[1578]  = A_iota[4][4][42];
    assign S_out[43]  = A_iota[0][0][43];
    assign S_out[107]  = A_iota[1][0][43];
    assign S_out[171]  = A_iota[2][0][43];
    assign S_out[235]  = A_iota[3][0][43];
    assign S_out[299]  = A_iota[4][0][43];
    assign S_out[363]  = A_iota[0][1][43];
    assign S_out[427]  = A_iota[1][1][43];
    assign S_out[491]  = A_iota[2][1][43];
    assign S_out[555]  = A_iota[3][1][43];
    assign S_out[619]  = A_iota[4][1][43];
    assign S_out[683]  = A_iota[0][2][43];
    assign S_out[747]  = A_iota[1][2][43];
    assign S_out[811]  = A_iota[2][2][43];
    assign S_out[875]  = A_iota[3][2][43];
    assign S_out[939]  = A_iota[4][2][43];
    assign S_out[1003]  = A_iota[0][3][43];
    assign S_out[1067]  = A_iota[1][3][43];
    assign S_out[1131]  = A_iota[2][3][43];
    assign S_out[1195]  = A_iota[3][3][43];
    assign S_out[1259]  = A_iota[4][3][43];
    assign S_out[1323]  = A_iota[0][4][43];
    assign S_out[1387]  = A_iota[1][4][43];
    assign S_out[1451]  = A_iota[2][4][43];
    assign S_out[1515]  = A_iota[3][4][43];
    assign S_out[1579]  = A_iota[4][4][43];
    assign S_out[44]  = A_iota[0][0][44];
    assign S_out[108]  = A_iota[1][0][44];
    assign S_out[172]  = A_iota[2][0][44];
    assign S_out[236]  = A_iota[3][0][44];
    assign S_out[300]  = A_iota[4][0][44];
    assign S_out[364]  = A_iota[0][1][44];
    assign S_out[428]  = A_iota[1][1][44];
    assign S_out[492]  = A_iota[2][1][44];
    assign S_out[556]  = A_iota[3][1][44];
    assign S_out[620]  = A_iota[4][1][44];
    assign S_out[684]  = A_iota[0][2][44];
    assign S_out[748]  = A_iota[1][2][44];
    assign S_out[812]  = A_iota[2][2][44];
    assign S_out[876]  = A_iota[3][2][44];
    assign S_out[940]  = A_iota[4][2][44];
    assign S_out[1004]  = A_iota[0][3][44];
    assign S_out[1068]  = A_iota[1][3][44];
    assign S_out[1132]  = A_iota[2][3][44];
    assign S_out[1196]  = A_iota[3][3][44];
    assign S_out[1260]  = A_iota[4][3][44];
    assign S_out[1324]  = A_iota[0][4][44];
    assign S_out[1388]  = A_iota[1][4][44];
    assign S_out[1452]  = A_iota[2][4][44];
    assign S_out[1516]  = A_iota[3][4][44];
    assign S_out[1580]  = A_iota[4][4][44];
    assign S_out[45]  = A_iota[0][0][45];
    assign S_out[109]  = A_iota[1][0][45];
    assign S_out[173]  = A_iota[2][0][45];
    assign S_out[237]  = A_iota[3][0][45];
    assign S_out[301]  = A_iota[4][0][45];
    assign S_out[365]  = A_iota[0][1][45];
    assign S_out[429]  = A_iota[1][1][45];
    assign S_out[493]  = A_iota[2][1][45];
    assign S_out[557]  = A_iota[3][1][45];
    assign S_out[621]  = A_iota[4][1][45];
    assign S_out[685]  = A_iota[0][2][45];
    assign S_out[749]  = A_iota[1][2][45];
    assign S_out[813]  = A_iota[2][2][45];
    assign S_out[877]  = A_iota[3][2][45];
    assign S_out[941]  = A_iota[4][2][45];
    assign S_out[1005]  = A_iota[0][3][45];
    assign S_out[1069]  = A_iota[1][3][45];
    assign S_out[1133]  = A_iota[2][3][45];
    assign S_out[1197]  = A_iota[3][3][45];
    assign S_out[1261]  = A_iota[4][3][45];
    assign S_out[1325]  = A_iota[0][4][45];
    assign S_out[1389]  = A_iota[1][4][45];
    assign S_out[1453]  = A_iota[2][4][45];
    assign S_out[1517]  = A_iota[3][4][45];
    assign S_out[1581]  = A_iota[4][4][45];
    assign S_out[46]  = A_iota[0][0][46];
    assign S_out[110]  = A_iota[1][0][46];
    assign S_out[174]  = A_iota[2][0][46];
    assign S_out[238]  = A_iota[3][0][46];
    assign S_out[302]  = A_iota[4][0][46];
    assign S_out[366]  = A_iota[0][1][46];
    assign S_out[430]  = A_iota[1][1][46];
    assign S_out[494]  = A_iota[2][1][46];
    assign S_out[558]  = A_iota[3][1][46];
    assign S_out[622]  = A_iota[4][1][46];
    assign S_out[686]  = A_iota[0][2][46];
    assign S_out[750]  = A_iota[1][2][46];
    assign S_out[814]  = A_iota[2][2][46];
    assign S_out[878]  = A_iota[3][2][46];
    assign S_out[942]  = A_iota[4][2][46];
    assign S_out[1006]  = A_iota[0][3][46];
    assign S_out[1070]  = A_iota[1][3][46];
    assign S_out[1134]  = A_iota[2][3][46];
    assign S_out[1198]  = A_iota[3][3][46];
    assign S_out[1262]  = A_iota[4][3][46];
    assign S_out[1326]  = A_iota[0][4][46];
    assign S_out[1390]  = A_iota[1][4][46];
    assign S_out[1454]  = A_iota[2][4][46];
    assign S_out[1518]  = A_iota[3][4][46];
    assign S_out[1582]  = A_iota[4][4][46];
    assign S_out[47]  = A_iota[0][0][47];
    assign S_out[111]  = A_iota[1][0][47];
    assign S_out[175]  = A_iota[2][0][47];
    assign S_out[239]  = A_iota[3][0][47];
    assign S_out[303]  = A_iota[4][0][47];
    assign S_out[367]  = A_iota[0][1][47];
    assign S_out[431]  = A_iota[1][1][47];
    assign S_out[495]  = A_iota[2][1][47];
    assign S_out[559]  = A_iota[3][1][47];
    assign S_out[623]  = A_iota[4][1][47];
    assign S_out[687]  = A_iota[0][2][47];
    assign S_out[751]  = A_iota[1][2][47];
    assign S_out[815]  = A_iota[2][2][47];
    assign S_out[879]  = A_iota[3][2][47];
    assign S_out[943]  = A_iota[4][2][47];
    assign S_out[1007]  = A_iota[0][3][47];
    assign S_out[1071]  = A_iota[1][3][47];
    assign S_out[1135]  = A_iota[2][3][47];
    assign S_out[1199]  = A_iota[3][3][47];
    assign S_out[1263]  = A_iota[4][3][47];
    assign S_out[1327]  = A_iota[0][4][47];
    assign S_out[1391]  = A_iota[1][4][47];
    assign S_out[1455]  = A_iota[2][4][47];
    assign S_out[1519]  = A_iota[3][4][47];
    assign S_out[1583]  = A_iota[4][4][47];
    assign S_out[48]  = A_iota[0][0][48];
    assign S_out[112]  = A_iota[1][0][48];
    assign S_out[176]  = A_iota[2][0][48];
    assign S_out[240]  = A_iota[3][0][48];
    assign S_out[304]  = A_iota[4][0][48];
    assign S_out[368]  = A_iota[0][1][48];
    assign S_out[432]  = A_iota[1][1][48];
    assign S_out[496]  = A_iota[2][1][48];
    assign S_out[560]  = A_iota[3][1][48];
    assign S_out[624]  = A_iota[4][1][48];
    assign S_out[688]  = A_iota[0][2][48];
    assign S_out[752]  = A_iota[1][2][48];
    assign S_out[816]  = A_iota[2][2][48];
    assign S_out[880]  = A_iota[3][2][48];
    assign S_out[944]  = A_iota[4][2][48];
    assign S_out[1008]  = A_iota[0][3][48];
    assign S_out[1072]  = A_iota[1][3][48];
    assign S_out[1136]  = A_iota[2][3][48];
    assign S_out[1200]  = A_iota[3][3][48];
    assign S_out[1264]  = A_iota[4][3][48];
    assign S_out[1328]  = A_iota[0][4][48];
    assign S_out[1392]  = A_iota[1][4][48];
    assign S_out[1456]  = A_iota[2][4][48];
    assign S_out[1520]  = A_iota[3][4][48];
    assign S_out[1584]  = A_iota[4][4][48];
    assign S_out[49]  = A_iota[0][0][49];
    assign S_out[113]  = A_iota[1][0][49];
    assign S_out[177]  = A_iota[2][0][49];
    assign S_out[241]  = A_iota[3][0][49];
    assign S_out[305]  = A_iota[4][0][49];
    assign S_out[369]  = A_iota[0][1][49];
    assign S_out[433]  = A_iota[1][1][49];
    assign S_out[497]  = A_iota[2][1][49];
    assign S_out[561]  = A_iota[3][1][49];
    assign S_out[625]  = A_iota[4][1][49];
    assign S_out[689]  = A_iota[0][2][49];
    assign S_out[753]  = A_iota[1][2][49];
    assign S_out[817]  = A_iota[2][2][49];
    assign S_out[881]  = A_iota[3][2][49];
    assign S_out[945]  = A_iota[4][2][49];
    assign S_out[1009]  = A_iota[0][3][49];
    assign S_out[1073]  = A_iota[1][3][49];
    assign S_out[1137]  = A_iota[2][3][49];
    assign S_out[1201]  = A_iota[3][3][49];
    assign S_out[1265]  = A_iota[4][3][49];
    assign S_out[1329]  = A_iota[0][4][49];
    assign S_out[1393]  = A_iota[1][4][49];
    assign S_out[1457]  = A_iota[2][4][49];
    assign S_out[1521]  = A_iota[3][4][49];
    assign S_out[1585]  = A_iota[4][4][49];
    assign S_out[50]  = A_iota[0][0][50];
    assign S_out[114]  = A_iota[1][0][50];
    assign S_out[178]  = A_iota[2][0][50];
    assign S_out[242]  = A_iota[3][0][50];
    assign S_out[306]  = A_iota[4][0][50];
    assign S_out[370]  = A_iota[0][1][50];
    assign S_out[434]  = A_iota[1][1][50];
    assign S_out[498]  = A_iota[2][1][50];
    assign S_out[562]  = A_iota[3][1][50];
    assign S_out[626]  = A_iota[4][1][50];
    assign S_out[690]  = A_iota[0][2][50];
    assign S_out[754]  = A_iota[1][2][50];
    assign S_out[818]  = A_iota[2][2][50];
    assign S_out[882]  = A_iota[3][2][50];
    assign S_out[946]  = A_iota[4][2][50];
    assign S_out[1010]  = A_iota[0][3][50];
    assign S_out[1074]  = A_iota[1][3][50];
    assign S_out[1138]  = A_iota[2][3][50];
    assign S_out[1202]  = A_iota[3][3][50];
    assign S_out[1266]  = A_iota[4][3][50];
    assign S_out[1330]  = A_iota[0][4][50];
    assign S_out[1394]  = A_iota[1][4][50];
    assign S_out[1458]  = A_iota[2][4][50];
    assign S_out[1522]  = A_iota[3][4][50];
    assign S_out[1586]  = A_iota[4][4][50];
    assign S_out[51]  = A_iota[0][0][51];
    assign S_out[115]  = A_iota[1][0][51];
    assign S_out[179]  = A_iota[2][0][51];
    assign S_out[243]  = A_iota[3][0][51];
    assign S_out[307]  = A_iota[4][0][51];
    assign S_out[371]  = A_iota[0][1][51];
    assign S_out[435]  = A_iota[1][1][51];
    assign S_out[499]  = A_iota[2][1][51];
    assign S_out[563]  = A_iota[3][1][51];
    assign S_out[627]  = A_iota[4][1][51];
    assign S_out[691]  = A_iota[0][2][51];
    assign S_out[755]  = A_iota[1][2][51];
    assign S_out[819]  = A_iota[2][2][51];
    assign S_out[883]  = A_iota[3][2][51];
    assign S_out[947]  = A_iota[4][2][51];
    assign S_out[1011]  = A_iota[0][3][51];
    assign S_out[1075]  = A_iota[1][3][51];
    assign S_out[1139]  = A_iota[2][3][51];
    assign S_out[1203]  = A_iota[3][3][51];
    assign S_out[1267]  = A_iota[4][3][51];
    assign S_out[1331]  = A_iota[0][4][51];
    assign S_out[1395]  = A_iota[1][4][51];
    assign S_out[1459]  = A_iota[2][4][51];
    assign S_out[1523]  = A_iota[3][4][51];
    assign S_out[1587]  = A_iota[4][4][51];
    assign S_out[52]  = A_iota[0][0][52];
    assign S_out[116]  = A_iota[1][0][52];
    assign S_out[180]  = A_iota[2][0][52];
    assign S_out[244]  = A_iota[3][0][52];
    assign S_out[308]  = A_iota[4][0][52];
    assign S_out[372]  = A_iota[0][1][52];
    assign S_out[436]  = A_iota[1][1][52];
    assign S_out[500]  = A_iota[2][1][52];
    assign S_out[564]  = A_iota[3][1][52];
    assign S_out[628]  = A_iota[4][1][52];
    assign S_out[692]  = A_iota[0][2][52];
    assign S_out[756]  = A_iota[1][2][52];
    assign S_out[820]  = A_iota[2][2][52];
    assign S_out[884]  = A_iota[3][2][52];
    assign S_out[948]  = A_iota[4][2][52];
    assign S_out[1012]  = A_iota[0][3][52];
    assign S_out[1076]  = A_iota[1][3][52];
    assign S_out[1140]  = A_iota[2][3][52];
    assign S_out[1204]  = A_iota[3][3][52];
    assign S_out[1268]  = A_iota[4][3][52];
    assign S_out[1332]  = A_iota[0][4][52];
    assign S_out[1396]  = A_iota[1][4][52];
    assign S_out[1460]  = A_iota[2][4][52];
    assign S_out[1524]  = A_iota[3][4][52];
    assign S_out[1588]  = A_iota[4][4][52];
    assign S_out[53]  = A_iota[0][0][53];
    assign S_out[117]  = A_iota[1][0][53];
    assign S_out[181]  = A_iota[2][0][53];
    assign S_out[245]  = A_iota[3][0][53];
    assign S_out[309]  = A_iota[4][0][53];
    assign S_out[373]  = A_iota[0][1][53];
    assign S_out[437]  = A_iota[1][1][53];
    assign S_out[501]  = A_iota[2][1][53];
    assign S_out[565]  = A_iota[3][1][53];
    assign S_out[629]  = A_iota[4][1][53];
    assign S_out[693]  = A_iota[0][2][53];
    assign S_out[757]  = A_iota[1][2][53];
    assign S_out[821]  = A_iota[2][2][53];
    assign S_out[885]  = A_iota[3][2][53];
    assign S_out[949]  = A_iota[4][2][53];
    assign S_out[1013]  = A_iota[0][3][53];
    assign S_out[1077]  = A_iota[1][3][53];
    assign S_out[1141]  = A_iota[2][3][53];
    assign S_out[1205]  = A_iota[3][3][53];
    assign S_out[1269]  = A_iota[4][3][53];
    assign S_out[1333]  = A_iota[0][4][53];
    assign S_out[1397]  = A_iota[1][4][53];
    assign S_out[1461]  = A_iota[2][4][53];
    assign S_out[1525]  = A_iota[3][4][53];
    assign S_out[1589]  = A_iota[4][4][53];
    assign S_out[54]  = A_iota[0][0][54];
    assign S_out[118]  = A_iota[1][0][54];
    assign S_out[182]  = A_iota[2][0][54];
    assign S_out[246]  = A_iota[3][0][54];
    assign S_out[310]  = A_iota[4][0][54];
    assign S_out[374]  = A_iota[0][1][54];
    assign S_out[438]  = A_iota[1][1][54];
    assign S_out[502]  = A_iota[2][1][54];
    assign S_out[566]  = A_iota[3][1][54];
    assign S_out[630]  = A_iota[4][1][54];
    assign S_out[694]  = A_iota[0][2][54];
    assign S_out[758]  = A_iota[1][2][54];
    assign S_out[822]  = A_iota[2][2][54];
    assign S_out[886]  = A_iota[3][2][54];
    assign S_out[950]  = A_iota[4][2][54];
    assign S_out[1014]  = A_iota[0][3][54];
    assign S_out[1078]  = A_iota[1][3][54];
    assign S_out[1142]  = A_iota[2][3][54];
    assign S_out[1206]  = A_iota[3][3][54];
    assign S_out[1270]  = A_iota[4][3][54];
    assign S_out[1334]  = A_iota[0][4][54];
    assign S_out[1398]  = A_iota[1][4][54];
    assign S_out[1462]  = A_iota[2][4][54];
    assign S_out[1526]  = A_iota[3][4][54];
    assign S_out[1590]  = A_iota[4][4][54];
    assign S_out[55]  = A_iota[0][0][55];
    assign S_out[119]  = A_iota[1][0][55];
    assign S_out[183]  = A_iota[2][0][55];
    assign S_out[247]  = A_iota[3][0][55];
    assign S_out[311]  = A_iota[4][0][55];
    assign S_out[375]  = A_iota[0][1][55];
    assign S_out[439]  = A_iota[1][1][55];
    assign S_out[503]  = A_iota[2][1][55];
    assign S_out[567]  = A_iota[3][1][55];
    assign S_out[631]  = A_iota[4][1][55];
    assign S_out[695]  = A_iota[0][2][55];
    assign S_out[759]  = A_iota[1][2][55];
    assign S_out[823]  = A_iota[2][2][55];
    assign S_out[887]  = A_iota[3][2][55];
    assign S_out[951]  = A_iota[4][2][55];
    assign S_out[1015]  = A_iota[0][3][55];
    assign S_out[1079]  = A_iota[1][3][55];
    assign S_out[1143]  = A_iota[2][3][55];
    assign S_out[1207]  = A_iota[3][3][55];
    assign S_out[1271]  = A_iota[4][3][55];
    assign S_out[1335]  = A_iota[0][4][55];
    assign S_out[1399]  = A_iota[1][4][55];
    assign S_out[1463]  = A_iota[2][4][55];
    assign S_out[1527]  = A_iota[3][4][55];
    assign S_out[1591]  = A_iota[4][4][55];
    assign S_out[56]  = A_iota[0][0][56];
    assign S_out[120]  = A_iota[1][0][56];
    assign S_out[184]  = A_iota[2][0][56];
    assign S_out[248]  = A_iota[3][0][56];
    assign S_out[312]  = A_iota[4][0][56];
    assign S_out[376]  = A_iota[0][1][56];
    assign S_out[440]  = A_iota[1][1][56];
    assign S_out[504]  = A_iota[2][1][56];
    assign S_out[568]  = A_iota[3][1][56];
    assign S_out[632]  = A_iota[4][1][56];
    assign S_out[696]  = A_iota[0][2][56];
    assign S_out[760]  = A_iota[1][2][56];
    assign S_out[824]  = A_iota[2][2][56];
    assign S_out[888]  = A_iota[3][2][56];
    assign S_out[952]  = A_iota[4][2][56];
    assign S_out[1016]  = A_iota[0][3][56];
    assign S_out[1080]  = A_iota[1][3][56];
    assign S_out[1144]  = A_iota[2][3][56];
    assign S_out[1208]  = A_iota[3][3][56];
    assign S_out[1272]  = A_iota[4][3][56];
    assign S_out[1336]  = A_iota[0][4][56];
    assign S_out[1400]  = A_iota[1][4][56];
    assign S_out[1464]  = A_iota[2][4][56];
    assign S_out[1528]  = A_iota[3][4][56];
    assign S_out[1592]  = A_iota[4][4][56];
    assign S_out[57]  = A_iota[0][0][57];
    assign S_out[121]  = A_iota[1][0][57];
    assign S_out[185]  = A_iota[2][0][57];
    assign S_out[249]  = A_iota[3][0][57];
    assign S_out[313]  = A_iota[4][0][57];
    assign S_out[377]  = A_iota[0][1][57];
    assign S_out[441]  = A_iota[1][1][57];
    assign S_out[505]  = A_iota[2][1][57];
    assign S_out[569]  = A_iota[3][1][57];
    assign S_out[633]  = A_iota[4][1][57];
    assign S_out[697]  = A_iota[0][2][57];
    assign S_out[761]  = A_iota[1][2][57];
    assign S_out[825]  = A_iota[2][2][57];
    assign S_out[889]  = A_iota[3][2][57];
    assign S_out[953]  = A_iota[4][2][57];
    assign S_out[1017]  = A_iota[0][3][57];
    assign S_out[1081]  = A_iota[1][3][57];
    assign S_out[1145]  = A_iota[2][3][57];
    assign S_out[1209]  = A_iota[3][3][57];
    assign S_out[1273]  = A_iota[4][3][57];
    assign S_out[1337]  = A_iota[0][4][57];
    assign S_out[1401]  = A_iota[1][4][57];
    assign S_out[1465]  = A_iota[2][4][57];
    assign S_out[1529]  = A_iota[3][4][57];
    assign S_out[1593]  = A_iota[4][4][57];
    assign S_out[58]  = A_iota[0][0][58];
    assign S_out[122]  = A_iota[1][0][58];
    assign S_out[186]  = A_iota[2][0][58];
    assign S_out[250]  = A_iota[3][0][58];
    assign S_out[314]  = A_iota[4][0][58];
    assign S_out[378]  = A_iota[0][1][58];
    assign S_out[442]  = A_iota[1][1][58];
    assign S_out[506]  = A_iota[2][1][58];
    assign S_out[570]  = A_iota[3][1][58];
    assign S_out[634]  = A_iota[4][1][58];
    assign S_out[698]  = A_iota[0][2][58];
    assign S_out[762]  = A_iota[1][2][58];
    assign S_out[826]  = A_iota[2][2][58];
    assign S_out[890]  = A_iota[3][2][58];
    assign S_out[954]  = A_iota[4][2][58];
    assign S_out[1018]  = A_iota[0][3][58];
    assign S_out[1082]  = A_iota[1][3][58];
    assign S_out[1146]  = A_iota[2][3][58];
    assign S_out[1210]  = A_iota[3][3][58];
    assign S_out[1274]  = A_iota[4][3][58];
    assign S_out[1338]  = A_iota[0][4][58];
    assign S_out[1402]  = A_iota[1][4][58];
    assign S_out[1466]  = A_iota[2][4][58];
    assign S_out[1530]  = A_iota[3][4][58];
    assign S_out[1594]  = A_iota[4][4][58];
    assign S_out[59]  = A_iota[0][0][59];
    assign S_out[123]  = A_iota[1][0][59];
    assign S_out[187]  = A_iota[2][0][59];
    assign S_out[251]  = A_iota[3][0][59];
    assign S_out[315]  = A_iota[4][0][59];
    assign S_out[379]  = A_iota[0][1][59];
    assign S_out[443]  = A_iota[1][1][59];
    assign S_out[507]  = A_iota[2][1][59];
    assign S_out[571]  = A_iota[3][1][59];
    assign S_out[635]  = A_iota[4][1][59];
    assign S_out[699]  = A_iota[0][2][59];
    assign S_out[763]  = A_iota[1][2][59];
    assign S_out[827]  = A_iota[2][2][59];
    assign S_out[891]  = A_iota[3][2][59];
    assign S_out[955]  = A_iota[4][2][59];
    assign S_out[1019]  = A_iota[0][3][59];
    assign S_out[1083]  = A_iota[1][3][59];
    assign S_out[1147]  = A_iota[2][3][59];
    assign S_out[1211]  = A_iota[3][3][59];
    assign S_out[1275]  = A_iota[4][3][59];
    assign S_out[1339]  = A_iota[0][4][59];
    assign S_out[1403]  = A_iota[1][4][59];
    assign S_out[1467]  = A_iota[2][4][59];
    assign S_out[1531]  = A_iota[3][4][59];
    assign S_out[1595]  = A_iota[4][4][59];
    assign S_out[60]  = A_iota[0][0][60];
    assign S_out[124]  = A_iota[1][0][60];
    assign S_out[188]  = A_iota[2][0][60];
    assign S_out[252]  = A_iota[3][0][60];
    assign S_out[316]  = A_iota[4][0][60];
    assign S_out[380]  = A_iota[0][1][60];
    assign S_out[444]  = A_iota[1][1][60];
    assign S_out[508]  = A_iota[2][1][60];
    assign S_out[572]  = A_iota[3][1][60];
    assign S_out[636]  = A_iota[4][1][60];
    assign S_out[700]  = A_iota[0][2][60];
    assign S_out[764]  = A_iota[1][2][60];
    assign S_out[828]  = A_iota[2][2][60];
    assign S_out[892]  = A_iota[3][2][60];
    assign S_out[956]  = A_iota[4][2][60];
    assign S_out[1020]  = A_iota[0][3][60];
    assign S_out[1084]  = A_iota[1][3][60];
    assign S_out[1148]  = A_iota[2][3][60];
    assign S_out[1212]  = A_iota[3][3][60];
    assign S_out[1276]  = A_iota[4][3][60];
    assign S_out[1340]  = A_iota[0][4][60];
    assign S_out[1404]  = A_iota[1][4][60];
    assign S_out[1468]  = A_iota[2][4][60];
    assign S_out[1532]  = A_iota[3][4][60];
    assign S_out[1596]  = A_iota[4][4][60];
    assign S_out[61]  = A_iota[0][0][61];
    assign S_out[125]  = A_iota[1][0][61];
    assign S_out[189]  = A_iota[2][0][61];
    assign S_out[253]  = A_iota[3][0][61];
    assign S_out[317]  = A_iota[4][0][61];
    assign S_out[381]  = A_iota[0][1][61];
    assign S_out[445]  = A_iota[1][1][61];
    assign S_out[509]  = A_iota[2][1][61];
    assign S_out[573]  = A_iota[3][1][61];
    assign S_out[637]  = A_iota[4][1][61];
    assign S_out[701]  = A_iota[0][2][61];
    assign S_out[765]  = A_iota[1][2][61];
    assign S_out[829]  = A_iota[2][2][61];
    assign S_out[893]  = A_iota[3][2][61];
    assign S_out[957]  = A_iota[4][2][61];
    assign S_out[1021]  = A_iota[0][3][61];
    assign S_out[1085]  = A_iota[1][3][61];
    assign S_out[1149]  = A_iota[2][3][61];
    assign S_out[1213]  = A_iota[3][3][61];
    assign S_out[1277]  = A_iota[4][3][61];
    assign S_out[1341]  = A_iota[0][4][61];
    assign S_out[1405]  = A_iota[1][4][61];
    assign S_out[1469]  = A_iota[2][4][61];
    assign S_out[1533]  = A_iota[3][4][61];
    assign S_out[1597]  = A_iota[4][4][61];
    assign S_out[62]  = A_iota[0][0][62];
    assign S_out[126]  = A_iota[1][0][62];
    assign S_out[190]  = A_iota[2][0][62];
    assign S_out[254]  = A_iota[3][0][62];
    assign S_out[318]  = A_iota[4][0][62];
    assign S_out[382]  = A_iota[0][1][62];
    assign S_out[446]  = A_iota[1][1][62];
    assign S_out[510]  = A_iota[2][1][62];
    assign S_out[574]  = A_iota[3][1][62];
    assign S_out[638]  = A_iota[4][1][62];
    assign S_out[702]  = A_iota[0][2][62];
    assign S_out[766]  = A_iota[1][2][62];
    assign S_out[830]  = A_iota[2][2][62];
    assign S_out[894]  = A_iota[3][2][62];
    assign S_out[958]  = A_iota[4][2][62];
    assign S_out[1022]  = A_iota[0][3][62];
    assign S_out[1086]  = A_iota[1][3][62];
    assign S_out[1150]  = A_iota[2][3][62];
    assign S_out[1214]  = A_iota[3][3][62];
    assign S_out[1278]  = A_iota[4][3][62];
    assign S_out[1342]  = A_iota[0][4][62];
    assign S_out[1406]  = A_iota[1][4][62];
    assign S_out[1470]  = A_iota[2][4][62];
    assign S_out[1534]  = A_iota[3][4][62];
    assign S_out[1598]  = A_iota[4][4][62];
    assign S_out[63]  = A_iota[0][0][63];
    assign S_out[127]  = A_iota[1][0][63];
    assign S_out[191]  = A_iota[2][0][63];
    assign S_out[255]  = A_iota[3][0][63];
    assign S_out[319]  = A_iota[4][0][63];
    assign S_out[383]  = A_iota[0][1][63];
    assign S_out[447]  = A_iota[1][1][63];
    assign S_out[511]  = A_iota[2][1][63];
    assign S_out[575]  = A_iota[3][1][63];
    assign S_out[639]  = A_iota[4][1][63];
    assign S_out[703]  = A_iota[0][2][63];
    assign S_out[767]  = A_iota[1][2][63];
    assign S_out[831]  = A_iota[2][2][63];
    assign S_out[895]  = A_iota[3][2][63];
    assign S_out[959]  = A_iota[4][2][63];
    assign S_out[1023]  = A_iota[0][3][63];
    assign S_out[1087]  = A_iota[1][3][63];
    assign S_out[1151]  = A_iota[2][3][63];
    assign S_out[1215]  = A_iota[3][3][63];
    assign S_out[1279]  = A_iota[4][3][63];
    assign S_out[1343]  = A_iota[0][4][63];
    assign S_out[1407]  = A_iota[1][4][63];
    assign S_out[1471]  = A_iota[2][4][63];
    assign S_out[1535]  = A_iota[3][4][63];
    assign S_out[1599]  = A_iota[4][4][63];
endmodule
